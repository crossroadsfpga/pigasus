`include "./src/struct_s.sv"
module non_fast_pattern_ht(clk,
    dout_0_0,dout_valid_0_0,
    dout_0_1,dout_valid_0_1,
    dout_0_2,dout_valid_0_2,
    dout_0_3,dout_valid_0_3,
    dout_0_4,dout_valid_0_4,
    dout_0_5,dout_valid_0_5,
    dout_0_6,dout_valid_0_6,
    dout_0_7,dout_valid_0_7,
    dout_0_8,dout_valid_0_8,
    dout_0_9,dout_valid_0_9,
    dout_0_10,dout_valid_0_10,
    dout_0_11,dout_valid_0_11,
    dout_0_12,dout_valid_0_12,
    dout_0_13,dout_valid_0_13,
    dout_0_14,dout_valid_0_14,
    dout_0_15,dout_valid_0_15,
    dout_1_0,dout_valid_1_0,
    dout_1_1,dout_valid_1_1,
    dout_1_2,dout_valid_1_2,
    dout_1_3,dout_valid_1_3,
    dout_1_4,dout_valid_1_4,
    dout_1_5,dout_valid_1_5,
    dout_1_6,dout_valid_1_6,
    dout_1_7,dout_valid_1_7,
    dout_1_8,dout_valid_1_8,
    dout_1_9,dout_valid_1_9,
    dout_1_10,dout_valid_1_10,
    dout_1_11,dout_valid_1_11,
    dout_1_12,dout_valid_1_12,
    dout_1_13,dout_valid_1_13,
    dout_1_14,dout_valid_1_14,
    dout_1_15,dout_valid_1_15,
    dout_2_0,dout_valid_2_0,
    dout_2_1,dout_valid_2_1,
    dout_2_2,dout_valid_2_2,
    dout_2_3,dout_valid_2_3,
    dout_2_4,dout_valid_2_4,
    dout_2_5,dout_valid_2_5,
    dout_2_6,dout_valid_2_6,
    dout_2_7,dout_valid_2_7,
    dout_2_8,dout_valid_2_8,
    dout_2_9,dout_valid_2_9,
    dout_2_10,dout_valid_2_10,
    dout_2_11,dout_valid_2_11,
    dout_2_12,dout_valid_2_12,
    dout_2_13,dout_valid_2_13,
    dout_2_14,dout_valid_2_14,
    dout_2_15,dout_valid_2_15,
    dout_3_0,dout_valid_3_0,
    dout_3_1,dout_valid_3_1,
    dout_3_2,dout_valid_3_2,
    dout_3_3,dout_valid_3_3,
    dout_3_4,dout_valid_3_4,
    dout_3_5,dout_valid_3_5,
    dout_3_6,dout_valid_3_6,
    dout_3_7,dout_valid_3_7,
    dout_3_8,dout_valid_3_8,
    dout_3_9,dout_valid_3_9,
    dout_3_10,dout_valid_3_10,
    dout_3_11,dout_valid_3_11,
    dout_3_12,dout_valid_3_12,
    dout_3_13,dout_valid_3_13,
    dout_3_14,dout_valid_3_14,
    dout_3_15,dout_valid_3_15,
    dout_4_0,dout_valid_4_0,
    dout_4_1,dout_valid_4_1,
    dout_4_2,dout_valid_4_2,
    dout_4_3,dout_valid_4_3,
    dout_4_4,dout_valid_4_4,
    dout_4_5,dout_valid_4_5,
    dout_4_6,dout_valid_4_6,
    dout_4_7,dout_valid_4_7,
    dout_4_8,dout_valid_4_8,
    dout_4_9,dout_valid_4_9,
    dout_4_10,dout_valid_4_10,
    dout_4_11,dout_valid_4_11,
    dout_4_12,dout_valid_4_12,
    dout_4_13,dout_valid_4_13,
    dout_4_14,dout_valid_4_14,
    dout_4_15,dout_valid_4_15,
    dout_5_0,dout_valid_5_0,
    dout_5_1,dout_valid_5_1,
    dout_5_2,dout_valid_5_2,
    dout_5_3,dout_valid_5_3,
    dout_5_4,dout_valid_5_4,
    dout_5_5,dout_valid_5_5,
    dout_5_6,dout_valid_5_6,
    dout_5_7,dout_valid_5_7,
    dout_5_8,dout_valid_5_8,
    dout_5_9,dout_valid_5_9,
    dout_5_10,dout_valid_5_10,
    dout_5_11,dout_valid_5_11,
    dout_5_12,dout_valid_5_12,
    dout_5_13,dout_valid_5_13,
    dout_5_14,dout_valid_5_14,
    dout_5_15,dout_valid_5_15,
    dout_6_0,dout_valid_6_0,
    dout_6_1,dout_valid_6_1,
    dout_6_2,dout_valid_6_2,
    dout_6_3,dout_valid_6_3,
    dout_6_4,dout_valid_6_4,
    dout_6_5,dout_valid_6_5,
    dout_6_6,dout_valid_6_6,
    dout_6_7,dout_valid_6_7,
    dout_6_8,dout_valid_6_8,
    dout_6_9,dout_valid_6_9,
    dout_6_10,dout_valid_6_10,
    dout_6_11,dout_valid_6_11,
    dout_6_12,dout_valid_6_12,
    dout_6_13,dout_valid_6_13,
    dout_6_14,dout_valid_6_14,
    dout_6_15,dout_valid_6_15,
    dout_7_0,dout_valid_7_0,
    dout_7_1,dout_valid_7_1,
    dout_7_2,dout_valid_7_2,
    dout_7_3,dout_valid_7_3,
    dout_7_4,dout_valid_7_4,
    dout_7_5,dout_valid_7_5,
    dout_7_6,dout_valid_7_6,
    dout_7_7,dout_valid_7_7,
    dout_7_8,dout_valid_7_8,
    dout_7_9,dout_valid_7_9,
    dout_7_10,dout_valid_7_10,
    dout_7_11,dout_valid_7_11,
    dout_7_12,dout_valid_7_12,
    dout_7_13,dout_valid_7_13,
    dout_7_14,dout_valid_7_14,
    dout_7_15,dout_valid_7_15,
    din,
    din_sop,
    din_valid
);

input clk;
input [NFP_DWIDTH-1:0] din;
input din_valid;
input din_sop;
output logic [NF_WIDTH-1:0] dout_0_0;
output logic dout_valid_0_0;
output logic [NF_WIDTH-1:0] dout_0_1;
output logic dout_valid_0_1;
output logic [NF_WIDTH-1:0] dout_0_2;
output logic dout_valid_0_2;
output logic [NF_WIDTH-1:0] dout_0_3;
output logic dout_valid_0_3;
output logic [NF_WIDTH-1:0] dout_0_4;
output logic dout_valid_0_4;
output logic [NF_WIDTH-1:0] dout_0_5;
output logic dout_valid_0_5;
output logic [NF_WIDTH-1:0] dout_0_6;
output logic dout_valid_0_6;
output logic [NF_WIDTH-1:0] dout_0_7;
output logic dout_valid_0_7;
output logic [NF_WIDTH-1:0] dout_0_8;
output logic dout_valid_0_8;
output logic [NF_WIDTH-1:0] dout_0_9;
output logic dout_valid_0_9;
output logic [NF_WIDTH-1:0] dout_0_10;
output logic dout_valid_0_10;
output logic [NF_WIDTH-1:0] dout_0_11;
output logic dout_valid_0_11;
output logic [NF_WIDTH-1:0] dout_0_12;
output logic dout_valid_0_12;
output logic [NF_WIDTH-1:0] dout_0_13;
output logic dout_valid_0_13;
output logic [NF_WIDTH-1:0] dout_0_14;
output logic dout_valid_0_14;
output logic [NF_WIDTH-1:0] dout_0_15;
output logic dout_valid_0_15;
output logic [NF_WIDTH-1:0] dout_1_0;
output logic dout_valid_1_0;
output logic [NF_WIDTH-1:0] dout_1_1;
output logic dout_valid_1_1;
output logic [NF_WIDTH-1:0] dout_1_2;
output logic dout_valid_1_2;
output logic [NF_WIDTH-1:0] dout_1_3;
output logic dout_valid_1_3;
output logic [NF_WIDTH-1:0] dout_1_4;
output logic dout_valid_1_4;
output logic [NF_WIDTH-1:0] dout_1_5;
output logic dout_valid_1_5;
output logic [NF_WIDTH-1:0] dout_1_6;
output logic dout_valid_1_6;
output logic [NF_WIDTH-1:0] dout_1_7;
output logic dout_valid_1_7;
output logic [NF_WIDTH-1:0] dout_1_8;
output logic dout_valid_1_8;
output logic [NF_WIDTH-1:0] dout_1_9;
output logic dout_valid_1_9;
output logic [NF_WIDTH-1:0] dout_1_10;
output logic dout_valid_1_10;
output logic [NF_WIDTH-1:0] dout_1_11;
output logic dout_valid_1_11;
output logic [NF_WIDTH-1:0] dout_1_12;
output logic dout_valid_1_12;
output logic [NF_WIDTH-1:0] dout_1_13;
output logic dout_valid_1_13;
output logic [NF_WIDTH-1:0] dout_1_14;
output logic dout_valid_1_14;
output logic [NF_WIDTH-1:0] dout_1_15;
output logic dout_valid_1_15;
output logic [NF_WIDTH-1:0] dout_2_0;
output logic dout_valid_2_0;
output logic [NF_WIDTH-1:0] dout_2_1;
output logic dout_valid_2_1;
output logic [NF_WIDTH-1:0] dout_2_2;
output logic dout_valid_2_2;
output logic [NF_WIDTH-1:0] dout_2_3;
output logic dout_valid_2_3;
output logic [NF_WIDTH-1:0] dout_2_4;
output logic dout_valid_2_4;
output logic [NF_WIDTH-1:0] dout_2_5;
output logic dout_valid_2_5;
output logic [NF_WIDTH-1:0] dout_2_6;
output logic dout_valid_2_6;
output logic [NF_WIDTH-1:0] dout_2_7;
output logic dout_valid_2_7;
output logic [NF_WIDTH-1:0] dout_2_8;
output logic dout_valid_2_8;
output logic [NF_WIDTH-1:0] dout_2_9;
output logic dout_valid_2_9;
output logic [NF_WIDTH-1:0] dout_2_10;
output logic dout_valid_2_10;
output logic [NF_WIDTH-1:0] dout_2_11;
output logic dout_valid_2_11;
output logic [NF_WIDTH-1:0] dout_2_12;
output logic dout_valid_2_12;
output logic [NF_WIDTH-1:0] dout_2_13;
output logic dout_valid_2_13;
output logic [NF_WIDTH-1:0] dout_2_14;
output logic dout_valid_2_14;
output logic [NF_WIDTH-1:0] dout_2_15;
output logic dout_valid_2_15;
output logic [NF_WIDTH-1:0] dout_3_0;
output logic dout_valid_3_0;
output logic [NF_WIDTH-1:0] dout_3_1;
output logic dout_valid_3_1;
output logic [NF_WIDTH-1:0] dout_3_2;
output logic dout_valid_3_2;
output logic [NF_WIDTH-1:0] dout_3_3;
output logic dout_valid_3_3;
output logic [NF_WIDTH-1:0] dout_3_4;
output logic dout_valid_3_4;
output logic [NF_WIDTH-1:0] dout_3_5;
output logic dout_valid_3_5;
output logic [NF_WIDTH-1:0] dout_3_6;
output logic dout_valid_3_6;
output logic [NF_WIDTH-1:0] dout_3_7;
output logic dout_valid_3_7;
output logic [NF_WIDTH-1:0] dout_3_8;
output logic dout_valid_3_8;
output logic [NF_WIDTH-1:0] dout_3_9;
output logic dout_valid_3_9;
output logic [NF_WIDTH-1:0] dout_3_10;
output logic dout_valid_3_10;
output logic [NF_WIDTH-1:0] dout_3_11;
output logic dout_valid_3_11;
output logic [NF_WIDTH-1:0] dout_3_12;
output logic dout_valid_3_12;
output logic [NF_WIDTH-1:0] dout_3_13;
output logic dout_valid_3_13;
output logic [NF_WIDTH-1:0] dout_3_14;
output logic dout_valid_3_14;
output logic [NF_WIDTH-1:0] dout_3_15;
output logic dout_valid_3_15;
output logic [NF_WIDTH-1:0] dout_4_0;
output logic dout_valid_4_0;
output logic [NF_WIDTH-1:0] dout_4_1;
output logic dout_valid_4_1;
output logic [NF_WIDTH-1:0] dout_4_2;
output logic dout_valid_4_2;
output logic [NF_WIDTH-1:0] dout_4_3;
output logic dout_valid_4_3;
output logic [NF_WIDTH-1:0] dout_4_4;
output logic dout_valid_4_4;
output logic [NF_WIDTH-1:0] dout_4_5;
output logic dout_valid_4_5;
output logic [NF_WIDTH-1:0] dout_4_6;
output logic dout_valid_4_6;
output logic [NF_WIDTH-1:0] dout_4_7;
output logic dout_valid_4_7;
output logic [NF_WIDTH-1:0] dout_4_8;
output logic dout_valid_4_8;
output logic [NF_WIDTH-1:0] dout_4_9;
output logic dout_valid_4_9;
output logic [NF_WIDTH-1:0] dout_4_10;
output logic dout_valid_4_10;
output logic [NF_WIDTH-1:0] dout_4_11;
output logic dout_valid_4_11;
output logic [NF_WIDTH-1:0] dout_4_12;
output logic dout_valid_4_12;
output logic [NF_WIDTH-1:0] dout_4_13;
output logic dout_valid_4_13;
output logic [NF_WIDTH-1:0] dout_4_14;
output logic dout_valid_4_14;
output logic [NF_WIDTH-1:0] dout_4_15;
output logic dout_valid_4_15;
output logic [NF_WIDTH-1:0] dout_5_0;
output logic dout_valid_5_0;
output logic [NF_WIDTH-1:0] dout_5_1;
output logic dout_valid_5_1;
output logic [NF_WIDTH-1:0] dout_5_2;
output logic dout_valid_5_2;
output logic [NF_WIDTH-1:0] dout_5_3;
output logic dout_valid_5_3;
output logic [NF_WIDTH-1:0] dout_5_4;
output logic dout_valid_5_4;
output logic [NF_WIDTH-1:0] dout_5_5;
output logic dout_valid_5_5;
output logic [NF_WIDTH-1:0] dout_5_6;
output logic dout_valid_5_6;
output logic [NF_WIDTH-1:0] dout_5_7;
output logic dout_valid_5_7;
output logic [NF_WIDTH-1:0] dout_5_8;
output logic dout_valid_5_8;
output logic [NF_WIDTH-1:0] dout_5_9;
output logic dout_valid_5_9;
output logic [NF_WIDTH-1:0] dout_5_10;
output logic dout_valid_5_10;
output logic [NF_WIDTH-1:0] dout_5_11;
output logic dout_valid_5_11;
output logic [NF_WIDTH-1:0] dout_5_12;
output logic dout_valid_5_12;
output logic [NF_WIDTH-1:0] dout_5_13;
output logic dout_valid_5_13;
output logic [NF_WIDTH-1:0] dout_5_14;
output logic dout_valid_5_14;
output logic [NF_WIDTH-1:0] dout_5_15;
output logic dout_valid_5_15;
output logic [NF_WIDTH-1:0] dout_6_0;
output logic dout_valid_6_0;
output logic [NF_WIDTH-1:0] dout_6_1;
output logic dout_valid_6_1;
output logic [NF_WIDTH-1:0] dout_6_2;
output logic dout_valid_6_2;
output logic [NF_WIDTH-1:0] dout_6_3;
output logic dout_valid_6_3;
output logic [NF_WIDTH-1:0] dout_6_4;
output logic dout_valid_6_4;
output logic [NF_WIDTH-1:0] dout_6_5;
output logic dout_valid_6_5;
output logic [NF_WIDTH-1:0] dout_6_6;
output logic dout_valid_6_6;
output logic [NF_WIDTH-1:0] dout_6_7;
output logic dout_valid_6_7;
output logic [NF_WIDTH-1:0] dout_6_8;
output logic dout_valid_6_8;
output logic [NF_WIDTH-1:0] dout_6_9;
output logic dout_valid_6_9;
output logic [NF_WIDTH-1:0] dout_6_10;
output logic dout_valid_6_10;
output logic [NF_WIDTH-1:0] dout_6_11;
output logic dout_valid_6_11;
output logic [NF_WIDTH-1:0] dout_6_12;
output logic dout_valid_6_12;
output logic [NF_WIDTH-1:0] dout_6_13;
output logic dout_valid_6_13;
output logic [NF_WIDTH-1:0] dout_6_14;
output logic dout_valid_6_14;
output logic [NF_WIDTH-1:0] dout_6_15;
output logic dout_valid_6_15;
output logic [NF_WIDTH-1:0] dout_7_0;
output logic dout_valid_7_0;
output logic [NF_WIDTH-1:0] dout_7_1;
output logic dout_valid_7_1;
output logic [NF_WIDTH-1:0] dout_7_2;
output logic dout_valid_7_2;
output logic [NF_WIDTH-1:0] dout_7_3;
output logic dout_valid_7_3;
output logic [NF_WIDTH-1:0] dout_7_4;
output logic dout_valid_7_4;
output logic [NF_WIDTH-1:0] dout_7_5;
output logic dout_valid_7_5;
output logic [NF_WIDTH-1:0] dout_7_6;
output logic dout_valid_7_6;
output logic [NF_WIDTH-1:0] dout_7_7;
output logic dout_valid_7_7;
output logic [NF_WIDTH-1:0] dout_7_8;
output logic dout_valid_7_8;
output logic [NF_WIDTH-1:0] dout_7_9;
output logic dout_valid_7_9;
output logic [NF_WIDTH-1:0] dout_7_10;
output logic dout_valid_7_10;
output logic [NF_WIDTH-1:0] dout_7_11;
output logic dout_valid_7_11;
output logic [NF_WIDTH-1:0] dout_7_12;
output logic dout_valid_7_12;
output logic [NF_WIDTH-1:0] dout_7_13;
output logic dout_valid_7_13;
output logic [NF_WIDTH-1:0] dout_7_14;
output logic dout_valid_7_14;
output logic [NF_WIDTH-1:0] dout_7_15;
output logic dout_valid_7_15;

reg  [17-1:0] addr_0_0;
logic din_valid_0_0;
wire addr_valid_0_0;
reg  [17-1:0] addr_0_1;
logic din_valid_0_1;
wire addr_valid_0_1;
reg  [17-1:0] addr_0_2;
logic din_valid_0_2;
wire addr_valid_0_2;
reg  [17-1:0] addr_0_3;
logic din_valid_0_3;
wire addr_valid_0_3;
reg  [17-1:0] addr_0_4;
logic din_valid_0_4;
wire addr_valid_0_4;
reg  [17-1:0] addr_0_5;
logic din_valid_0_5;
wire addr_valid_0_5;
reg  [17-1:0] addr_0_6;
logic din_valid_0_6;
wire addr_valid_0_6;
reg  [17-1:0] addr_0_7;
logic din_valid_0_7;
wire addr_valid_0_7;
reg  [17-1:0] addr_0_8;
logic din_valid_0_8;
wire addr_valid_0_8;
reg  [17-1:0] addr_0_9;
logic din_valid_0_9;
wire addr_valid_0_9;
reg  [17-1:0] addr_0_10;
logic din_valid_0_10;
wire addr_valid_0_10;
reg  [17-1:0] addr_0_11;
logic din_valid_0_11;
wire addr_valid_0_11;
reg  [17-1:0] addr_0_12;
logic din_valid_0_12;
wire addr_valid_0_12;
reg  [17-1:0] addr_0_13;
logic din_valid_0_13;
wire addr_valid_0_13;
reg  [17-1:0] addr_0_14;
logic din_valid_0_14;
wire addr_valid_0_14;
reg  [17-1:0] addr_0_15;
logic din_valid_0_15;
wire addr_valid_0_15;
reg  [13-1:0] addr_1_0;
logic din_valid_1_0;
wire addr_valid_1_0;
reg  [13-1:0] addr_1_1;
logic din_valid_1_1;
wire addr_valid_1_1;
reg  [13-1:0] addr_1_2;
logic din_valid_1_2;
wire addr_valid_1_2;
reg  [13-1:0] addr_1_3;
logic din_valid_1_3;
wire addr_valid_1_3;
reg  [13-1:0] addr_1_4;
logic din_valid_1_4;
wire addr_valid_1_4;
reg  [13-1:0] addr_1_5;
logic din_valid_1_5;
wire addr_valid_1_5;
reg  [13-1:0] addr_1_6;
logic din_valid_1_6;
wire addr_valid_1_6;
reg  [13-1:0] addr_1_7;
logic din_valid_1_7;
wire addr_valid_1_7;
reg  [13-1:0] addr_1_8;
logic din_valid_1_8;
wire addr_valid_1_8;
reg  [13-1:0] addr_1_9;
logic din_valid_1_9;
wire addr_valid_1_9;
reg  [13-1:0] addr_1_10;
logic din_valid_1_10;
wire addr_valid_1_10;
reg  [13-1:0] addr_1_11;
logic din_valid_1_11;
wire addr_valid_1_11;
reg  [13-1:0] addr_1_12;
logic din_valid_1_12;
wire addr_valid_1_12;
reg  [13-1:0] addr_1_13;
logic din_valid_1_13;
wire addr_valid_1_13;
reg  [13-1:0] addr_1_14;
logic din_valid_1_14;
wire addr_valid_1_14;
reg  [13-1:0] addr_1_15;
logic din_valid_1_15;
wire addr_valid_1_15;
reg  [13-1:0] addr_2_0;
logic din_valid_2_0;
wire addr_valid_2_0;
reg  [13-1:0] addr_2_1;
logic din_valid_2_1;
wire addr_valid_2_1;
reg  [13-1:0] addr_2_2;
logic din_valid_2_2;
wire addr_valid_2_2;
reg  [13-1:0] addr_2_3;
logic din_valid_2_3;
wire addr_valid_2_3;
reg  [13-1:0] addr_2_4;
logic din_valid_2_4;
wire addr_valid_2_4;
reg  [13-1:0] addr_2_5;
logic din_valid_2_5;
wire addr_valid_2_5;
reg  [13-1:0] addr_2_6;
logic din_valid_2_6;
wire addr_valid_2_6;
reg  [13-1:0] addr_2_7;
logic din_valid_2_7;
wire addr_valid_2_7;
reg  [13-1:0] addr_2_8;
logic din_valid_2_8;
wire addr_valid_2_8;
reg  [13-1:0] addr_2_9;
logic din_valid_2_9;
wire addr_valid_2_9;
reg  [13-1:0] addr_2_10;
logic din_valid_2_10;
wire addr_valid_2_10;
reg  [13-1:0] addr_2_11;
logic din_valid_2_11;
wire addr_valid_2_11;
reg  [13-1:0] addr_2_12;
logic din_valid_2_12;
wire addr_valid_2_12;
reg  [13-1:0] addr_2_13;
logic din_valid_2_13;
wire addr_valid_2_13;
reg  [13-1:0] addr_2_14;
logic din_valid_2_14;
wire addr_valid_2_14;
reg  [13-1:0] addr_2_15;
logic din_valid_2_15;
wire addr_valid_2_15;
reg  [13-1:0] addr_3_0;
logic din_valid_3_0;
wire addr_valid_3_0;
reg  [13-1:0] addr_3_1;
logic din_valid_3_1;
wire addr_valid_3_1;
reg  [13-1:0] addr_3_2;
logic din_valid_3_2;
wire addr_valid_3_2;
reg  [13-1:0] addr_3_3;
logic din_valid_3_3;
wire addr_valid_3_3;
reg  [13-1:0] addr_3_4;
logic din_valid_3_4;
wire addr_valid_3_4;
reg  [13-1:0] addr_3_5;
logic din_valid_3_5;
wire addr_valid_3_5;
reg  [13-1:0] addr_3_6;
logic din_valid_3_6;
wire addr_valid_3_6;
reg  [13-1:0] addr_3_7;
logic din_valid_3_7;
wire addr_valid_3_7;
reg  [13-1:0] addr_3_8;
logic din_valid_3_8;
wire addr_valid_3_8;
reg  [13-1:0] addr_3_9;
logic din_valid_3_9;
wire addr_valid_3_9;
reg  [13-1:0] addr_3_10;
logic din_valid_3_10;
wire addr_valid_3_10;
reg  [13-1:0] addr_3_11;
logic din_valid_3_11;
wire addr_valid_3_11;
reg  [13-1:0] addr_3_12;
logic din_valid_3_12;
wire addr_valid_3_12;
reg  [13-1:0] addr_3_13;
logic din_valid_3_13;
wire addr_valid_3_13;
reg  [13-1:0] addr_3_14;
logic din_valid_3_14;
wire addr_valid_3_14;
reg  [13-1:0] addr_3_15;
logic din_valid_3_15;
wire addr_valid_3_15;
reg  [13-1:0] addr_4_0;
logic din_valid_4_0;
wire addr_valid_4_0;
reg  [13-1:0] addr_4_1;
logic din_valid_4_1;
wire addr_valid_4_1;
reg  [13-1:0] addr_4_2;
logic din_valid_4_2;
wire addr_valid_4_2;
reg  [13-1:0] addr_4_3;
logic din_valid_4_3;
wire addr_valid_4_3;
reg  [13-1:0] addr_4_4;
logic din_valid_4_4;
wire addr_valid_4_4;
reg  [13-1:0] addr_4_5;
logic din_valid_4_5;
wire addr_valid_4_5;
reg  [13-1:0] addr_4_6;
logic din_valid_4_6;
wire addr_valid_4_6;
reg  [13-1:0] addr_4_7;
logic din_valid_4_7;
wire addr_valid_4_7;
reg  [13-1:0] addr_4_8;
logic din_valid_4_8;
wire addr_valid_4_8;
reg  [13-1:0] addr_4_9;
logic din_valid_4_9;
wire addr_valid_4_9;
reg  [13-1:0] addr_4_10;
logic din_valid_4_10;
wire addr_valid_4_10;
reg  [13-1:0] addr_4_11;
logic din_valid_4_11;
wire addr_valid_4_11;
reg  [13-1:0] addr_4_12;
logic din_valid_4_12;
wire addr_valid_4_12;
reg  [13-1:0] addr_4_13;
logic din_valid_4_13;
wire addr_valid_4_13;
reg  [13-1:0] addr_4_14;
logic din_valid_4_14;
wire addr_valid_4_14;
reg  [13-1:0] addr_4_15;
logic din_valid_4_15;
wire addr_valid_4_15;
reg  [12-1:0] addr_5_0;
logic din_valid_5_0;
wire addr_valid_5_0;
reg  [12-1:0] addr_5_1;
logic din_valid_5_1;
wire addr_valid_5_1;
reg  [12-1:0] addr_5_2;
logic din_valid_5_2;
wire addr_valid_5_2;
reg  [12-1:0] addr_5_3;
logic din_valid_5_3;
wire addr_valid_5_3;
reg  [12-1:0] addr_5_4;
logic din_valid_5_4;
wire addr_valid_5_4;
reg  [12-1:0] addr_5_5;
logic din_valid_5_5;
wire addr_valid_5_5;
reg  [12-1:0] addr_5_6;
logic din_valid_5_6;
wire addr_valid_5_6;
reg  [12-1:0] addr_5_7;
logic din_valid_5_7;
wire addr_valid_5_7;
reg  [12-1:0] addr_5_8;
logic din_valid_5_8;
wire addr_valid_5_8;
reg  [12-1:0] addr_5_9;
logic din_valid_5_9;
wire addr_valid_5_9;
reg  [12-1:0] addr_5_10;
logic din_valid_5_10;
wire addr_valid_5_10;
reg  [12-1:0] addr_5_11;
logic din_valid_5_11;
wire addr_valid_5_11;
reg  [12-1:0] addr_5_12;
logic din_valid_5_12;
wire addr_valid_5_12;
reg  [12-1:0] addr_5_13;
logic din_valid_5_13;
wire addr_valid_5_13;
reg  [12-1:0] addr_5_14;
logic din_valid_5_14;
wire addr_valid_5_14;
reg  [12-1:0] addr_5_15;
logic din_valid_5_15;
wire addr_valid_5_15;
reg  [11-1:0] addr_6_0;
logic din_valid_6_0;
wire addr_valid_6_0;
reg  [11-1:0] addr_6_1;
logic din_valid_6_1;
wire addr_valid_6_1;
reg  [11-1:0] addr_6_2;
logic din_valid_6_2;
wire addr_valid_6_2;
reg  [11-1:0] addr_6_3;
logic din_valid_6_3;
wire addr_valid_6_3;
reg  [11-1:0] addr_6_4;
logic din_valid_6_4;
wire addr_valid_6_4;
reg  [11-1:0] addr_6_5;
logic din_valid_6_5;
wire addr_valid_6_5;
reg  [11-1:0] addr_6_6;
logic din_valid_6_6;
wire addr_valid_6_6;
reg  [11-1:0] addr_6_7;
logic din_valid_6_7;
wire addr_valid_6_7;
reg  [11-1:0] addr_6_8;
logic din_valid_6_8;
wire addr_valid_6_8;
reg  [11-1:0] addr_6_9;
logic din_valid_6_9;
wire addr_valid_6_9;
reg  [11-1:0] addr_6_10;
logic din_valid_6_10;
wire addr_valid_6_10;
reg  [11-1:0] addr_6_11;
logic din_valid_6_11;
wire addr_valid_6_11;
reg  [11-1:0] addr_6_12;
logic din_valid_6_12;
wire addr_valid_6_12;
reg  [11-1:0] addr_6_13;
logic din_valid_6_13;
wire addr_valid_6_13;
reg  [11-1:0] addr_6_14;
logic din_valid_6_14;
wire addr_valid_6_14;
reg  [11-1:0] addr_6_15;
logic din_valid_6_15;
wire addr_valid_6_15;
reg  [10-1:0] addr_7_0;
logic din_valid_7_0;
wire addr_valid_7_0;
reg  [10-1:0] addr_7_1;
logic din_valid_7_1;
wire addr_valid_7_1;
reg  [10-1:0] addr_7_2;
logic din_valid_7_2;
wire addr_valid_7_2;
reg  [10-1:0] addr_7_3;
logic din_valid_7_3;
wire addr_valid_7_3;
reg  [10-1:0] addr_7_4;
logic din_valid_7_4;
wire addr_valid_7_4;
reg  [10-1:0] addr_7_5;
logic din_valid_7_5;
wire addr_valid_7_5;
reg  [10-1:0] addr_7_6;
logic din_valid_7_6;
wire addr_valid_7_6;
reg  [10-1:0] addr_7_7;
logic din_valid_7_7;
wire addr_valid_7_7;
reg  [10-1:0] addr_7_8;
logic din_valid_7_8;
wire addr_valid_7_8;
reg  [10-1:0] addr_7_9;
logic din_valid_7_9;
wire addr_valid_7_9;
reg  [10-1:0] addr_7_10;
logic din_valid_7_10;
wire addr_valid_7_10;
reg  [10-1:0] addr_7_11;
logic din_valid_7_11;
wire addr_valid_7_11;
reg  [10-1:0] addr_7_12;
logic din_valid_7_12;
wire addr_valid_7_12;
reg  [10-1:0] addr_7_13;
logic din_valid_7_13;
wire addr_valid_7_13;
reg  [10-1:0] addr_7_14;
logic din_valid_7_14;
wire addr_valid_7_14;
reg  [10-1:0] addr_7_15;
logic din_valid_7_15;
wire addr_valid_7_15;

logic din_valid_reg;
logic [63:0] din_reg;

// Doing all necessary multiplies per input byte
wire [(16+7)*8-1:0] padded_din;

wire [23:0] din_0_ab0;
wire [23:0] din_0_ab1;
wire [23:0] din_0_ab2;
wire [23:0] din_0_ab3;
wire [23:0] din_1_ab0;
wire [23:0] din_1_ab1;
wire [23:0] din_1_ab2;
wire [23:0] din_1_ab3;
wire [23:0] din_2_ab0;
wire [23:0] din_2_ab1;
wire [23:0] din_2_ab2;
wire [23:0] din_2_ab3;
wire [23:0] din_3_ab0;
wire [23:0] din_3_ab1;
wire [23:0] din_3_ab2;
wire [23:0] din_3_ab3;
wire [23:0] din_4_ab0;
wire [23:0] din_4_ab1;
wire [23:0] din_4_ab2;
wire [23:0] din_4_ab3;
wire [23:0] din_5_ab0;
wire [23:0] din_5_ab1;
wire [23:0] din_5_ab2;
wire [23:0] din_5_ab3;
wire [23:0] din_6_ab0;
wire [23:0] din_6_ab1;
wire [23:0] din_6_ab2;
wire [23:0] din_6_ab3;
wire [23:0] din_7_ab0;
wire [23:0] din_7_ab1;
wire [23:0] din_7_ab2;
wire [23:0] din_7_ab3;
wire [23:0] din_8_ab0;
wire [23:0] din_8_ab1;
wire [23:0] din_8_ab2;
wire [23:0] din_8_ab3;
wire [23:0] din_9_ab0;
wire [23:0] din_9_ab1;
wire [23:0] din_9_ab2;
wire [23:0] din_9_ab3;
wire [23:0] din_10_ab0;
wire [23:0] din_10_ab1;
wire [23:0] din_10_ab2;
wire [23:0] din_10_ab3;
wire [23:0] din_11_ab0;
wire [23:0] din_11_ab1;
wire [23:0] din_11_ab2;
wire [23:0] din_11_ab3;
wire [23:0] din_12_ab0;
wire [23:0] din_12_ab1;
wire [23:0] din_12_ab2;
wire [23:0] din_12_ab3;
wire [23:0] din_13_ab0;
wire [23:0] din_13_ab1;
wire [23:0] din_13_ab2;
wire [23:0] din_13_ab3;
wire [23:0] din_14_ab0;
wire [23:0] din_14_ab1;
wire [23:0] din_14_ab2;
wire [23:0] din_14_ab3;
wire [23:0] din_15_ab0;
wire [23:0] din_15_ab1;
wire [23:0] din_15_ab2;
wire [23:0] din_15_ab3;
wire [23:0] din_16_ab0;
wire [23:0] din_16_ab1;
wire [23:0] din_16_ab2;
wire [23:0] din_16_ab3;
wire [23:0] din_17_ab0;
wire [23:0] din_17_ab1;
wire [23:0] din_17_ab2;
wire [23:0] din_17_ab3;
wire [23:0] din_18_ab0;
wire [23:0] din_18_ab1;
wire [23:0] din_18_ab2;
wire [23:0] din_18_ab3;
wire [23:0] din_19_ab0;
wire [23:0] din_19_ab1;
wire [23:0] din_19_ab2;
wire [23:0] din_19_ab3;
wire [23:0] din_20_ab0;
wire [23:0] din_20_ab1;
wire [23:0] din_20_ab2;
wire [23:0] din_20_ab3;
wire [23:0] din_21_ab0;
wire [23:0] din_21_ab1;
wire [23:0] din_21_ab2;
wire [23:0] din_21_ab3;
wire [23:0] din_22_ab0;
wire [23:0] din_22_ab1;
wire [23:0] din_22_ab2;
wire [23:0] din_22_ab3;

assign padded_din = {din[16*8-1:0], din_reg[63:8]};

mul_hash din_0_mul_hash (
    .clk(clk),
    .a(padded_din[0*8+:8]), 
    .ab0(din_0_ab0),                 
    .ab1(din_0_ab1), 
    .ab2(din_0_ab2),                 
    .ab3(din_0_ab3)
);

mul_hash din_1_mul_hash (
    .clk(clk),
    .a(padded_din[1*8+:8]), 
    .ab0(din_1_ab0),                 
    .ab1(din_1_ab1), 
    .ab2(din_1_ab2),                 
    .ab3(din_1_ab3)
);

mul_hash din_2_mul_hash (
    .clk(clk),
    .a(padded_din[2*8+:8]), 
    .ab0(din_2_ab0),                 
    .ab1(din_2_ab1), 
    .ab2(din_2_ab2),                 
    .ab3(din_2_ab3)
);

mul_hash din_3_mul_hash (
    .clk(clk),
    .a(padded_din[3*8+:8]), 
    .ab0(din_3_ab0),                 
    .ab1(din_3_ab1), 
    .ab2(din_3_ab2),                 
    .ab3(din_3_ab3)
);

mul_hash din_4_mul_hash (
    .clk(clk),
    .a(padded_din[4*8+:8]), 
    .ab0(din_4_ab0),                 
    .ab1(din_4_ab1), 
    .ab2(din_4_ab2),                 
    .ab3(din_4_ab3)
);

mul_hash din_5_mul_hash (
    .clk(clk),
    .a(padded_din[5*8+:8]), 
    .ab0(din_5_ab0),                 
    .ab1(din_5_ab1), 
    .ab2(din_5_ab2),                 
    .ab3(din_5_ab3)
);

mul_hash din_6_mul_hash (
    .clk(clk),
    .a(padded_din[6*8+:8]), 
    .ab0(din_6_ab0),                 
    .ab1(din_6_ab1), 
    .ab2(din_6_ab2),                 
    .ab3(din_6_ab3)
);

mul_hash din_7_mul_hash (
    .clk(clk),
    .a(padded_din[7*8+:8]), 
    .ab0(din_7_ab0),                 
    .ab1(din_7_ab1), 
    .ab2(din_7_ab2),                 
    .ab3(din_7_ab3)
);

mul_hash din_8_mul_hash (
    .clk(clk),
    .a(padded_din[8*8+:8]), 
    .ab0(din_8_ab0),                 
    .ab1(din_8_ab1), 
    .ab2(din_8_ab2),                 
    .ab3(din_8_ab3)
);

mul_hash din_9_mul_hash (
    .clk(clk),
    .a(padded_din[9*8+:8]), 
    .ab0(din_9_ab0),                 
    .ab1(din_9_ab1), 
    .ab2(din_9_ab2),                 
    .ab3(din_9_ab3)
);

mul_hash din_10_mul_hash (
    .clk(clk),
    .a(padded_din[10*8+:8]), 
    .ab0(din_10_ab0),                 
    .ab1(din_10_ab1), 
    .ab2(din_10_ab2),                 
    .ab3(din_10_ab3)
);

mul_hash din_11_mul_hash (
    .clk(clk),
    .a(padded_din[11*8+:8]), 
    .ab0(din_11_ab0),                 
    .ab1(din_11_ab1), 
    .ab2(din_11_ab2),                 
    .ab3(din_11_ab3)
);

mul_hash din_12_mul_hash (
    .clk(clk),
    .a(padded_din[12*8+:8]), 
    .ab0(din_12_ab0),                 
    .ab1(din_12_ab1), 
    .ab2(din_12_ab2),                 
    .ab3(din_12_ab3)
);

mul_hash din_13_mul_hash (
    .clk(clk),
    .a(padded_din[13*8+:8]), 
    .ab0(din_13_ab0),                 
    .ab1(din_13_ab1), 
    .ab2(din_13_ab2),                 
    .ab3(din_13_ab3)
);

mul_hash din_14_mul_hash (
    .clk(clk),
    .a(padded_din[14*8+:8]), 
    .ab0(din_14_ab0),                 
    .ab1(din_14_ab1), 
    .ab2(din_14_ab2),                 
    .ab3(din_14_ab3)
);

mul_hash din_15_mul_hash (
    .clk(clk),
    .a(padded_din[15*8+:8]), 
    .ab0(din_15_ab0),                 
    .ab1(din_15_ab1), 
    .ab2(din_15_ab2),                 
    .ab3(din_15_ab3)
);

mul_hash din_16_mul_hash (
    .clk(clk),
    .a(padded_din[16*8+:8]), 
    .ab0(din_16_ab0),                 
    .ab1(din_16_ab1), 
    .ab2(din_16_ab2),                 
    .ab3(din_16_ab3)
);

mul_hash din_17_mul_hash (
    .clk(clk),
    .a(padded_din[17*8+:8]), 
    .ab0(din_17_ab0),                 
    .ab1(din_17_ab1), 
    .ab2(din_17_ab2),                 
    .ab3(din_17_ab3)
);

mul_hash din_18_mul_hash (
    .clk(clk),
    .a(padded_din[18*8+:8]), 
    .ab0(din_18_ab0),                 
    .ab1(din_18_ab1), 
    .ab2(din_18_ab2),                 
    .ab3(din_18_ab3)
);

mul_hash din_19_mul_hash (
    .clk(clk),
    .a(padded_din[19*8+:8]), 
    .ab0(din_19_ab0),                 
    .ab1(din_19_ab1), 
    .ab2(din_19_ab2),                 
    .ab3(din_19_ab3)
);

mul_hash din_20_mul_hash (
    .clk(clk),
    .a(padded_din[20*8+:8]), 
    .ab0(din_20_ab0),                 
    .ab1(din_20_ab1), 
    .ab2(din_20_ab2),                 
    .ab3(din_20_ab3)
);

mul_hash din_21_mul_hash (
    .clk(clk),
    .a(padded_din[21*8+:8]), 
    .ab0(din_21_ab0),                 
    .ab1(din_21_ab1), 
    .ab2(din_21_ab2),                 
    .ab3(din_21_ab3)
);

mul_hash din_22_mul_hash (
    .clk(clk),
    .a(padded_din[22*8+:8]), 
    .ab0(din_22_ab0),                 
    .ab1(din_22_ab1), 
    .ab2(din_22_ab2),                 
    .ab3(din_22_ab3)
);



//Valid signals
assign din_valid_0_0 = din_valid & din_valid_reg;
assign din_valid_0_1 = din_valid & din_valid_reg;
assign din_valid_0_2 = din_valid & din_valid_reg;
assign din_valid_0_3 = din_valid & din_valid_reg;
assign din_valid_0_4 = din_valid & din_valid_reg;
assign din_valid_0_5 = din_valid & din_valid_reg;
assign din_valid_0_6 = din_valid & din_valid_reg;
assign din_valid_0_7 = din_valid;
assign din_valid_0_8 = din_valid;
assign din_valid_0_9 = din_valid;
assign din_valid_0_10 = din_valid;
assign din_valid_0_11 = din_valid;
assign din_valid_0_12 = din_valid;
assign din_valid_0_13 = din_valid;
assign din_valid_0_14 = din_valid;
assign din_valid_0_15 = din_valid;

assign din_valid_1_0 = din_valid & din_valid_reg;
assign din_valid_1_1 = din_valid & din_valid_reg;
assign din_valid_1_2 = din_valid & din_valid_reg;
assign din_valid_1_3 = din_valid & din_valid_reg;
assign din_valid_1_4 = din_valid & din_valid_reg;
assign din_valid_1_5 = din_valid & din_valid_reg;
assign din_valid_1_6 = din_valid;
assign din_valid_1_7 = din_valid;
assign din_valid_1_8 = din_valid;
assign din_valid_1_9 = din_valid;
assign din_valid_1_10 = din_valid;
assign din_valid_1_11 = din_valid;
assign din_valid_1_12 = din_valid;
assign din_valid_1_13 = din_valid;
assign din_valid_1_14 = din_valid;
assign din_valid_1_15 = din_valid;

assign din_valid_2_0 = din_valid & din_valid_reg;
assign din_valid_2_1 = din_valid & din_valid_reg;
assign din_valid_2_2 = din_valid & din_valid_reg;
assign din_valid_2_3 = din_valid & din_valid_reg;
assign din_valid_2_4 = din_valid & din_valid_reg;
assign din_valid_2_5 = din_valid;
assign din_valid_2_6 = din_valid;
assign din_valid_2_7 = din_valid;
assign din_valid_2_8 = din_valid;
assign din_valid_2_9 = din_valid;
assign din_valid_2_10 = din_valid;
assign din_valid_2_11 = din_valid;
assign din_valid_2_12 = din_valid;
assign din_valid_2_13 = din_valid;
assign din_valid_2_14 = din_valid;
assign din_valid_2_15 = din_valid;

assign din_valid_3_0 = din_valid & din_valid_reg;
assign din_valid_3_1 = din_valid & din_valid_reg;
assign din_valid_3_2 = din_valid & din_valid_reg;
assign din_valid_3_3 = din_valid & din_valid_reg;
assign din_valid_3_4 = din_valid;
assign din_valid_3_5 = din_valid;
assign din_valid_3_6 = din_valid;
assign din_valid_3_7 = din_valid;
assign din_valid_3_8 = din_valid;
assign din_valid_3_9 = din_valid;
assign din_valid_3_10 = din_valid;
assign din_valid_3_11 = din_valid;
assign din_valid_3_12 = din_valid;
assign din_valid_3_13 = din_valid;
assign din_valid_3_14 = din_valid;
assign din_valid_3_15 = din_valid;

assign din_valid_4_0 = din_valid & din_valid_reg;
assign din_valid_4_1 = din_valid & din_valid_reg;
assign din_valid_4_2 = din_valid & din_valid_reg;
assign din_valid_4_3 = din_valid;
assign din_valid_4_4 = din_valid;
assign din_valid_4_5 = din_valid;
assign din_valid_4_6 = din_valid;
assign din_valid_4_7 = din_valid;
assign din_valid_4_8 = din_valid;
assign din_valid_4_9 = din_valid;
assign din_valid_4_10 = din_valid;
assign din_valid_4_11 = din_valid;
assign din_valid_4_12 = din_valid;
assign din_valid_4_13 = din_valid;
assign din_valid_4_14 = din_valid;
assign din_valid_4_15 = din_valid;

assign din_valid_5_0 = din_valid & din_valid_reg;
assign din_valid_5_1 = din_valid & din_valid_reg;
assign din_valid_5_2 = din_valid;
assign din_valid_5_3 = din_valid;
assign din_valid_5_4 = din_valid;
assign din_valid_5_5 = din_valid;
assign din_valid_5_6 = din_valid;
assign din_valid_5_7 = din_valid;
assign din_valid_5_8 = din_valid;
assign din_valid_5_9 = din_valid;
assign din_valid_5_10 = din_valid;
assign din_valid_5_11 = din_valid;
assign din_valid_5_12 = din_valid;
assign din_valid_5_13 = din_valid;
assign din_valid_5_14 = din_valid;
assign din_valid_5_15 = din_valid;

assign din_valid_6_0 = din_valid & din_valid_reg;
assign din_valid_6_1 = din_valid;
assign din_valid_6_2 = din_valid;
assign din_valid_6_3 = din_valid;
assign din_valid_6_4 = din_valid;
assign din_valid_6_5 = din_valid;
assign din_valid_6_6 = din_valid;
assign din_valid_6_7 = din_valid;
assign din_valid_6_8 = din_valid;
assign din_valid_6_9 = din_valid;
assign din_valid_6_10 = din_valid;
assign din_valid_6_11 = din_valid;
assign din_valid_6_12 = din_valid;
assign din_valid_6_13 = din_valid;
assign din_valid_6_14 = din_valid;
assign din_valid_6_15 = din_valid;

assign din_valid_7_0 = din_valid;
assign din_valid_7_1 = din_valid;
assign din_valid_7_2 = din_valid;
assign din_valid_7_3 = din_valid;
assign din_valid_7_4 = din_valid;
assign din_valid_7_5 = din_valid;
assign din_valid_7_6 = din_valid;
assign din_valid_7_7 = din_valid;
assign din_valid_7_8 = din_valid;
assign din_valid_7_9 = din_valid;
assign din_valid_7_10 = din_valid;
assign din_valid_7_11 = din_valid;
assign din_valid_7_12 = din_valid;
assign din_valid_7_13 = din_valid;
assign din_valid_7_14 = din_valid;
assign din_valid_7_15 = din_valid;


always @ (posedge clk) begin
    din_reg <= din[NFP_DWIDTH-1:NFP_DWIDTH-64];
    din_valid_reg <= din_valid;
end

// 12 cycles latency for valid signals
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_0_pipe (
    .clk(clk),.din(din_valid_0_0),.dout(addr_valid_0_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_1_pipe (
    .clk(clk),.din(din_valid_0_1),.dout(addr_valid_0_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_2_pipe (
    .clk(clk),.din(din_valid_0_2),.dout(addr_valid_0_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_3_pipe (
    .clk(clk),.din(din_valid_0_3),.dout(addr_valid_0_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_4_pipe (
    .clk(clk),.din(din_valid_0_4),.dout(addr_valid_0_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_5_pipe (
    .clk(clk),.din(din_valid_0_5),.dout(addr_valid_0_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_6_pipe (
    .clk(clk),.din(din_valid_0_6),.dout(addr_valid_0_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_7_pipe (
    .clk(clk),.din(din_valid_0_7),.dout(addr_valid_0_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_8_pipe (
    .clk(clk),.din(din_valid_0_8),.dout(addr_valid_0_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_9_pipe (
    .clk(clk),.din(din_valid_0_9),.dout(addr_valid_0_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_10_pipe (
    .clk(clk),.din(din_valid_0_10),.dout(addr_valid_0_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_11_pipe (
    .clk(clk),.din(din_valid_0_11),.dout(addr_valid_0_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_12_pipe (
    .clk(clk),.din(din_valid_0_12),.dout(addr_valid_0_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_13_pipe (
    .clk(clk),.din(din_valid_0_13),.dout(addr_valid_0_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_14_pipe (
    .clk(clk),.din(din_valid_0_14),.dout(addr_valid_0_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_0_15_pipe (
    .clk(clk),.din(din_valid_0_15),.dout(addr_valid_0_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_0_pipe (
    .clk(clk),.din(din_valid_1_0),.dout(addr_valid_1_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_1_pipe (
    .clk(clk),.din(din_valid_1_1),.dout(addr_valid_1_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_2_pipe (
    .clk(clk),.din(din_valid_1_2),.dout(addr_valid_1_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_3_pipe (
    .clk(clk),.din(din_valid_1_3),.dout(addr_valid_1_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_4_pipe (
    .clk(clk),.din(din_valid_1_4),.dout(addr_valid_1_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_5_pipe (
    .clk(clk),.din(din_valid_1_5),.dout(addr_valid_1_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_6_pipe (
    .clk(clk),.din(din_valid_1_6),.dout(addr_valid_1_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_7_pipe (
    .clk(clk),.din(din_valid_1_7),.dout(addr_valid_1_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_8_pipe (
    .clk(clk),.din(din_valid_1_8),.dout(addr_valid_1_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_9_pipe (
    .clk(clk),.din(din_valid_1_9),.dout(addr_valid_1_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_10_pipe (
    .clk(clk),.din(din_valid_1_10),.dout(addr_valid_1_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_11_pipe (
    .clk(clk),.din(din_valid_1_11),.dout(addr_valid_1_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_12_pipe (
    .clk(clk),.din(din_valid_1_12),.dout(addr_valid_1_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_13_pipe (
    .clk(clk),.din(din_valid_1_13),.dout(addr_valid_1_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_14_pipe (
    .clk(clk),.din(din_valid_1_14),.dout(addr_valid_1_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_1_15_pipe (
    .clk(clk),.din(din_valid_1_15),.dout(addr_valid_1_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_0_pipe (
    .clk(clk),.din(din_valid_2_0),.dout(addr_valid_2_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_1_pipe (
    .clk(clk),.din(din_valid_2_1),.dout(addr_valid_2_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_2_pipe (
    .clk(clk),.din(din_valid_2_2),.dout(addr_valid_2_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_3_pipe (
    .clk(clk),.din(din_valid_2_3),.dout(addr_valid_2_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_4_pipe (
    .clk(clk),.din(din_valid_2_4),.dout(addr_valid_2_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_5_pipe (
    .clk(clk),.din(din_valid_2_5),.dout(addr_valid_2_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_6_pipe (
    .clk(clk),.din(din_valid_2_6),.dout(addr_valid_2_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_7_pipe (
    .clk(clk),.din(din_valid_2_7),.dout(addr_valid_2_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_8_pipe (
    .clk(clk),.din(din_valid_2_8),.dout(addr_valid_2_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_9_pipe (
    .clk(clk),.din(din_valid_2_9),.dout(addr_valid_2_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_10_pipe (
    .clk(clk),.din(din_valid_2_10),.dout(addr_valid_2_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_11_pipe (
    .clk(clk),.din(din_valid_2_11),.dout(addr_valid_2_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_12_pipe (
    .clk(clk),.din(din_valid_2_12),.dout(addr_valid_2_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_13_pipe (
    .clk(clk),.din(din_valid_2_13),.dout(addr_valid_2_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_14_pipe (
    .clk(clk),.din(din_valid_2_14),.dout(addr_valid_2_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_2_15_pipe (
    .clk(clk),.din(din_valid_2_15),.dout(addr_valid_2_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_0_pipe (
    .clk(clk),.din(din_valid_3_0),.dout(addr_valid_3_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_1_pipe (
    .clk(clk),.din(din_valid_3_1),.dout(addr_valid_3_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_2_pipe (
    .clk(clk),.din(din_valid_3_2),.dout(addr_valid_3_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_3_pipe (
    .clk(clk),.din(din_valid_3_3),.dout(addr_valid_3_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_4_pipe (
    .clk(clk),.din(din_valid_3_4),.dout(addr_valid_3_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_5_pipe (
    .clk(clk),.din(din_valid_3_5),.dout(addr_valid_3_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_6_pipe (
    .clk(clk),.din(din_valid_3_6),.dout(addr_valid_3_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_7_pipe (
    .clk(clk),.din(din_valid_3_7),.dout(addr_valid_3_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_8_pipe (
    .clk(clk),.din(din_valid_3_8),.dout(addr_valid_3_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_9_pipe (
    .clk(clk),.din(din_valid_3_9),.dout(addr_valid_3_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_10_pipe (
    .clk(clk),.din(din_valid_3_10),.dout(addr_valid_3_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_11_pipe (
    .clk(clk),.din(din_valid_3_11),.dout(addr_valid_3_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_12_pipe (
    .clk(clk),.din(din_valid_3_12),.dout(addr_valid_3_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_13_pipe (
    .clk(clk),.din(din_valid_3_13),.dout(addr_valid_3_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_14_pipe (
    .clk(clk),.din(din_valid_3_14),.dout(addr_valid_3_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_3_15_pipe (
    .clk(clk),.din(din_valid_3_15),.dout(addr_valid_3_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_0_pipe (
    .clk(clk),.din(din_valid_4_0),.dout(addr_valid_4_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_1_pipe (
    .clk(clk),.din(din_valid_4_1),.dout(addr_valid_4_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_2_pipe (
    .clk(clk),.din(din_valid_4_2),.dout(addr_valid_4_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_3_pipe (
    .clk(clk),.din(din_valid_4_3),.dout(addr_valid_4_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_4_pipe (
    .clk(clk),.din(din_valid_4_4),.dout(addr_valid_4_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_5_pipe (
    .clk(clk),.din(din_valid_4_5),.dout(addr_valid_4_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_6_pipe (
    .clk(clk),.din(din_valid_4_6),.dout(addr_valid_4_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_7_pipe (
    .clk(clk),.din(din_valid_4_7),.dout(addr_valid_4_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_8_pipe (
    .clk(clk),.din(din_valid_4_8),.dout(addr_valid_4_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_9_pipe (
    .clk(clk),.din(din_valid_4_9),.dout(addr_valid_4_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_10_pipe (
    .clk(clk),.din(din_valid_4_10),.dout(addr_valid_4_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_11_pipe (
    .clk(clk),.din(din_valid_4_11),.dout(addr_valid_4_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_12_pipe (
    .clk(clk),.din(din_valid_4_12),.dout(addr_valid_4_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_13_pipe (
    .clk(clk),.din(din_valid_4_13),.dout(addr_valid_4_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_14_pipe (
    .clk(clk),.din(din_valid_4_14),.dout(addr_valid_4_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_4_15_pipe (
    .clk(clk),.din(din_valid_4_15),.dout(addr_valid_4_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_0_pipe (
    .clk(clk),.din(din_valid_5_0),.dout(addr_valid_5_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_1_pipe (
    .clk(clk),.din(din_valid_5_1),.dout(addr_valid_5_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_2_pipe (
    .clk(clk),.din(din_valid_5_2),.dout(addr_valid_5_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_3_pipe (
    .clk(clk),.din(din_valid_5_3),.dout(addr_valid_5_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_4_pipe (
    .clk(clk),.din(din_valid_5_4),.dout(addr_valid_5_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_5_pipe (
    .clk(clk),.din(din_valid_5_5),.dout(addr_valid_5_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_6_pipe (
    .clk(clk),.din(din_valid_5_6),.dout(addr_valid_5_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_7_pipe (
    .clk(clk),.din(din_valid_5_7),.dout(addr_valid_5_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_8_pipe (
    .clk(clk),.din(din_valid_5_8),.dout(addr_valid_5_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_9_pipe (
    .clk(clk),.din(din_valid_5_9),.dout(addr_valid_5_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_10_pipe (
    .clk(clk),.din(din_valid_5_10),.dout(addr_valid_5_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_11_pipe (
    .clk(clk),.din(din_valid_5_11),.dout(addr_valid_5_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_12_pipe (
    .clk(clk),.din(din_valid_5_12),.dout(addr_valid_5_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_13_pipe (
    .clk(clk),.din(din_valid_5_13),.dout(addr_valid_5_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_14_pipe (
    .clk(clk),.din(din_valid_5_14),.dout(addr_valid_5_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_5_15_pipe (
    .clk(clk),.din(din_valid_5_15),.dout(addr_valid_5_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_0_pipe (
    .clk(clk),.din(din_valid_6_0),.dout(addr_valid_6_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_1_pipe (
    .clk(clk),.din(din_valid_6_1),.dout(addr_valid_6_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_2_pipe (
    .clk(clk),.din(din_valid_6_2),.dout(addr_valid_6_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_3_pipe (
    .clk(clk),.din(din_valid_6_3),.dout(addr_valid_6_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_4_pipe (
    .clk(clk),.din(din_valid_6_4),.dout(addr_valid_6_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_5_pipe (
    .clk(clk),.din(din_valid_6_5),.dout(addr_valid_6_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_6_pipe (
    .clk(clk),.din(din_valid_6_6),.dout(addr_valid_6_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_7_pipe (
    .clk(clk),.din(din_valid_6_7),.dout(addr_valid_6_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_8_pipe (
    .clk(clk),.din(din_valid_6_8),.dout(addr_valid_6_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_9_pipe (
    .clk(clk),.din(din_valid_6_9),.dout(addr_valid_6_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_10_pipe (
    .clk(clk),.din(din_valid_6_10),.dout(addr_valid_6_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_11_pipe (
    .clk(clk),.din(din_valid_6_11),.dout(addr_valid_6_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_12_pipe (
    .clk(clk),.din(din_valid_6_12),.dout(addr_valid_6_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_13_pipe (
    .clk(clk),.din(din_valid_6_13),.dout(addr_valid_6_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_14_pipe (
    .clk(clk),.din(din_valid_6_14),.dout(addr_valid_6_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_6_15_pipe (
    .clk(clk),.din(din_valid_6_15),.dout(addr_valid_6_15));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_0_pipe (
    .clk(clk),.din(din_valid_7_0),.dout(addr_valid_7_0));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_1_pipe (
    .clk(clk),.din(din_valid_7_1),.dout(addr_valid_7_1));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_2_pipe (
    .clk(clk),.din(din_valid_7_2),.dout(addr_valid_7_2));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_3_pipe (
    .clk(clk),.din(din_valid_7_3),.dout(addr_valid_7_3));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_4_pipe (
    .clk(clk),.din(din_valid_7_4),.dout(addr_valid_7_4));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_5_pipe (
    .clk(clk),.din(din_valid_7_5),.dout(addr_valid_7_5));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_6_pipe (
    .clk(clk),.din(din_valid_7_6),.dout(addr_valid_7_6));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_7_pipe (
    .clk(clk),.din(din_valid_7_7),.dout(addr_valid_7_7));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_8_pipe (
    .clk(clk),.din(din_valid_7_8),.dout(addr_valid_7_8));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_9_pipe (
    .clk(clk),.din(din_valid_7_9),.dout(addr_valid_7_9));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_10_pipe (
    .clk(clk),.din(din_valid_7_10),.dout(addr_valid_7_10));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_11_pipe (
    .clk(clk),.din(din_valid_7_11),.dout(addr_valid_7_11));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_12_pipe (
    .clk(clk),.din(din_valid_7_12),.dout(addr_valid_7_12));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_13_pipe (
    .clk(clk),.din(din_valid_7_13),.dout(addr_valid_7_13));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_14_pipe (
    .clk(clk),.din(din_valid_7_14),.dout(addr_valid_7_14));
hyper_pipe #(.NUM_PIPES(12)) addr_valid_7_15_pipe (
    .clk(clk),.din(din_valid_7_15),.dout(addr_valid_7_15));

// Multiply accumulation step. 
// Mask and Nbits is dependent on bucket number
// data selection is dependent on first byte location
acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_0_calc (
  .clk(clk), .p(addr_0_0),
  .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
  .a1b0(din_1_ab0), .a1b1(din_1_ab1), .a1b2(din_1_ab2), .a1b3(din_1_ab3),
  .a2b0(din_2_ab0), .a2b1(din_2_ab1), .a2b2(din_2_ab2),
  .a3b0(din_3_ab0), .a3b1(din_3_ab1), .a3b2(din_3_ab2),
  .a4b0(din_4_ab0), .a4b1(din_4_ab1),
  .a5b0(din_5_ab0), .a5b1(din_5_ab1),
  .a6b0(din_6_ab0),
  .a7b0(din_7_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_1_calc (
  .clk(clk), .p(addr_0_1),
  .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
  .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2), .a1b3(din_2_ab3),
  .a2b0(din_3_ab0), .a2b1(din_3_ab1), .a2b2(din_3_ab2),
  .a3b0(din_4_ab0), .a3b1(din_4_ab1), .a3b2(din_4_ab2),
  .a4b0(din_5_ab0), .a4b1(din_5_ab1),
  .a5b0(din_6_ab0), .a5b1(din_6_ab1),
  .a6b0(din_7_ab0),
  .a7b0(din_8_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_2_calc (
  .clk(clk), .p(addr_0_2),
  .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
  .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2), .a1b3(din_3_ab3),
  .a2b0(din_4_ab0), .a2b1(din_4_ab1), .a2b2(din_4_ab2),
  .a3b0(din_5_ab0), .a3b1(din_5_ab1), .a3b2(din_5_ab2),
  .a4b0(din_6_ab0), .a4b1(din_6_ab1),
  .a5b0(din_7_ab0), .a5b1(din_7_ab1),
  .a6b0(din_8_ab0),
  .a7b0(din_9_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_3_calc (
  .clk(clk), .p(addr_0_3),
  .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
  .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2), .a1b3(din_4_ab3),
  .a2b0(din_5_ab0), .a2b1(din_5_ab1), .a2b2(din_5_ab2),
  .a3b0(din_6_ab0), .a3b1(din_6_ab1), .a3b2(din_6_ab2),
  .a4b0(din_7_ab0), .a4b1(din_7_ab1),
  .a5b0(din_8_ab0), .a5b1(din_8_ab1),
  .a6b0(din_9_ab0),
  .a7b0(din_10_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_4_calc (
  .clk(clk), .p(addr_0_4),
  .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
  .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2), .a1b3(din_5_ab3),
  .a2b0(din_6_ab0), .a2b1(din_6_ab1), .a2b2(din_6_ab2),
  .a3b0(din_7_ab0), .a3b1(din_7_ab1), .a3b2(din_7_ab2),
  .a4b0(din_8_ab0), .a4b1(din_8_ab1),
  .a5b0(din_9_ab0), .a5b1(din_9_ab1),
  .a6b0(din_10_ab0),
  .a7b0(din_11_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_5_calc (
  .clk(clk), .p(addr_0_5),
  .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
  .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2), .a1b3(din_6_ab3),
  .a2b0(din_7_ab0), .a2b1(din_7_ab1), .a2b2(din_7_ab2),
  .a3b0(din_8_ab0), .a3b1(din_8_ab1), .a3b2(din_8_ab2),
  .a4b0(din_9_ab0), .a4b1(din_9_ab1),
  .a5b0(din_10_ab0), .a5b1(din_10_ab1),
  .a6b0(din_11_ab0),
  .a7b0(din_12_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_6_calc (
  .clk(clk), .p(addr_0_6),
  .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
  .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2), .a1b3(din_7_ab3),
  .a2b0(din_8_ab0), .a2b1(din_8_ab1), .a2b2(din_8_ab2),
  .a3b0(din_9_ab0), .a3b1(din_9_ab1), .a3b2(din_9_ab2),
  .a4b0(din_10_ab0), .a4b1(din_10_ab1),
  .a5b0(din_11_ab0), .a5b1(din_11_ab1),
  .a6b0(din_12_ab0),
  .a7b0(din_13_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_7_calc (
  .clk(clk), .p(addr_0_7),
  .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
  .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2), .a1b3(din_8_ab3),
  .a2b0(din_9_ab0), .a2b1(din_9_ab1), .a2b2(din_9_ab2),
  .a3b0(din_10_ab0), .a3b1(din_10_ab1), .a3b2(din_10_ab2),
  .a4b0(din_11_ab0), .a4b1(din_11_ab1),
  .a5b0(din_12_ab0), .a5b1(din_12_ab1),
  .a6b0(din_13_ab0),
  .a7b0(din_14_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_8_calc (
  .clk(clk), .p(addr_0_8),
  .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
  .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2), .a1b3(din_9_ab3),
  .a2b0(din_10_ab0), .a2b1(din_10_ab1), .a2b2(din_10_ab2),
  .a3b0(din_11_ab0), .a3b1(din_11_ab1), .a3b2(din_11_ab2),
  .a4b0(din_12_ab0), .a4b1(din_12_ab1),
  .a5b0(din_13_ab0), .a5b1(din_13_ab1),
  .a6b0(din_14_ab0),
  .a7b0(din_15_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_9_calc (
  .clk(clk), .p(addr_0_9),
  .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
  .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2), .a1b3(din_10_ab3),
  .a2b0(din_11_ab0), .a2b1(din_11_ab1), .a2b2(din_11_ab2),
  .a3b0(din_12_ab0), .a3b1(din_12_ab1), .a3b2(din_12_ab2),
  .a4b0(din_13_ab0), .a4b1(din_13_ab1),
  .a5b0(din_14_ab0), .a5b1(din_14_ab1),
  .a6b0(din_15_ab0),
  .a7b0(din_16_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_10_calc (
  .clk(clk), .p(addr_0_10),
  .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
  .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2), .a1b3(din_11_ab3),
  .a2b0(din_12_ab0), .a2b1(din_12_ab1), .a2b2(din_12_ab2),
  .a3b0(din_13_ab0), .a3b1(din_13_ab1), .a3b2(din_13_ab2),
  .a4b0(din_14_ab0), .a4b1(din_14_ab1),
  .a5b0(din_15_ab0), .a5b1(din_15_ab1),
  .a6b0(din_16_ab0),
  .a7b0(din_17_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_11_calc (
  .clk(clk), .p(addr_0_11),
  .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
  .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2), .a1b3(din_12_ab3),
  .a2b0(din_13_ab0), .a2b1(din_13_ab1), .a2b2(din_13_ab2),
  .a3b0(din_14_ab0), .a3b1(din_14_ab1), .a3b2(din_14_ab2),
  .a4b0(din_15_ab0), .a4b1(din_15_ab1),
  .a5b0(din_16_ab0), .a5b1(din_16_ab1),
  .a6b0(din_17_ab0),
  .a7b0(din_18_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_12_calc (
  .clk(clk), .p(addr_0_12),
  .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
  .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2), .a1b3(din_13_ab3),
  .a2b0(din_14_ab0), .a2b1(din_14_ab1), .a2b2(din_14_ab2),
  .a3b0(din_15_ab0), .a3b1(din_15_ab1), .a3b2(din_15_ab2),
  .a4b0(din_16_ab0), .a4b1(din_16_ab1),
  .a5b0(din_17_ab0), .a5b1(din_17_ab1),
  .a6b0(din_18_ab0),
  .a7b0(din_19_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_13_calc (
  .clk(clk), .p(addr_0_13),
  .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
  .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2), .a1b3(din_14_ab3),
  .a2b0(din_15_ab0), .a2b1(din_15_ab1), .a2b2(din_15_ab2),
  .a3b0(din_16_ab0), .a3b1(din_16_ab1), .a3b2(din_16_ab2),
  .a4b0(din_17_ab0), .a4b1(din_17_ab1),
  .a5b0(din_18_ab0), .a5b1(din_18_ab1),
  .a6b0(din_19_ab0),
  .a7b0(din_20_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_14_calc (
  .clk(clk), .p(addr_0_14),
  .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
  .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2), .a1b3(din_15_ab3),
  .a2b0(din_16_ab0), .a2b1(din_16_ab1), .a2b2(din_16_ab2),
  .a3b0(din_17_ab0), .a3b1(din_17_ab1), .a3b2(din_17_ab2),
  .a4b0(din_18_ab0), .a4b1(din_18_ab1),
  .a5b0(din_19_ab0), .a5b1(din_19_ab1),
  .a6b0(din_20_ab0),
  .a7b0(din_21_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(17)
) addr_0_15_calc (
  .clk(clk), .p(addr_0_15),
  .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
  .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2), .a1b3(din_16_ab3),
  .a2b0(din_17_ab0), .a2b1(din_17_ab1), .a2b2(din_17_ab2),
  .a3b0(din_18_ab0), .a3b1(din_18_ab1), .a3b2(din_18_ab2),
  .a4b0(din_19_ab0), .a4b1(din_19_ab1),
  .a5b0(din_20_ab0), .a5b1(din_20_ab1),
  .a6b0(din_21_ab0),
  .a7b0(din_22_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_0_calc (
  .clk(clk), .p(addr_1_0),
  .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
  .a1b0(din_1_ab0), .a1b1(din_1_ab1), .a1b2(din_1_ab2), .a1b3(din_1_ab3),
  .a2b0(din_2_ab0), .a2b1(din_2_ab1), .a2b2(din_2_ab2),
  .a3b0(din_3_ab0), .a3b1(din_3_ab1), .a3b2(din_3_ab2),
  .a4b0(din_4_ab0), .a4b1(din_4_ab1),
  .a5b0(din_5_ab0), .a5b1(din_5_ab1),
  .a6b0(din_6_ab0),
  .a7b0(din_7_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_1_calc (
  .clk(clk), .p(addr_1_1),
  .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
  .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2), .a1b3(din_2_ab3),
  .a2b0(din_3_ab0), .a2b1(din_3_ab1), .a2b2(din_3_ab2),
  .a3b0(din_4_ab0), .a3b1(din_4_ab1), .a3b2(din_4_ab2),
  .a4b0(din_5_ab0), .a4b1(din_5_ab1),
  .a5b0(din_6_ab0), .a5b1(din_6_ab1),
  .a6b0(din_7_ab0),
  .a7b0(din_8_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_2_calc (
  .clk(clk), .p(addr_1_2),
  .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
  .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2), .a1b3(din_3_ab3),
  .a2b0(din_4_ab0), .a2b1(din_4_ab1), .a2b2(din_4_ab2),
  .a3b0(din_5_ab0), .a3b1(din_5_ab1), .a3b2(din_5_ab2),
  .a4b0(din_6_ab0), .a4b1(din_6_ab1),
  .a5b0(din_7_ab0), .a5b1(din_7_ab1),
  .a6b0(din_8_ab0),
  .a7b0(din_9_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_3_calc (
  .clk(clk), .p(addr_1_3),
  .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
  .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2), .a1b3(din_4_ab3),
  .a2b0(din_5_ab0), .a2b1(din_5_ab1), .a2b2(din_5_ab2),
  .a3b0(din_6_ab0), .a3b1(din_6_ab1), .a3b2(din_6_ab2),
  .a4b0(din_7_ab0), .a4b1(din_7_ab1),
  .a5b0(din_8_ab0), .a5b1(din_8_ab1),
  .a6b0(din_9_ab0),
  .a7b0(din_10_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_4_calc (
  .clk(clk), .p(addr_1_4),
  .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
  .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2), .a1b3(din_5_ab3),
  .a2b0(din_6_ab0), .a2b1(din_6_ab1), .a2b2(din_6_ab2),
  .a3b0(din_7_ab0), .a3b1(din_7_ab1), .a3b2(din_7_ab2),
  .a4b0(din_8_ab0), .a4b1(din_8_ab1),
  .a5b0(din_9_ab0), .a5b1(din_9_ab1),
  .a6b0(din_10_ab0),
  .a7b0(din_11_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_5_calc (
  .clk(clk), .p(addr_1_5),
  .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
  .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2), .a1b3(din_6_ab3),
  .a2b0(din_7_ab0), .a2b1(din_7_ab1), .a2b2(din_7_ab2),
  .a3b0(din_8_ab0), .a3b1(din_8_ab1), .a3b2(din_8_ab2),
  .a4b0(din_9_ab0), .a4b1(din_9_ab1),
  .a5b0(din_10_ab0), .a5b1(din_10_ab1),
  .a6b0(din_11_ab0),
  .a7b0(din_12_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_6_calc (
  .clk(clk), .p(addr_1_6),
  .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
  .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2), .a1b3(din_7_ab3),
  .a2b0(din_8_ab0), .a2b1(din_8_ab1), .a2b2(din_8_ab2),
  .a3b0(din_9_ab0), .a3b1(din_9_ab1), .a3b2(din_9_ab2),
  .a4b0(din_10_ab0), .a4b1(din_10_ab1),
  .a5b0(din_11_ab0), .a5b1(din_11_ab1),
  .a6b0(din_12_ab0),
  .a7b0(din_13_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_7_calc (
  .clk(clk), .p(addr_1_7),
  .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
  .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2), .a1b3(din_8_ab3),
  .a2b0(din_9_ab0), .a2b1(din_9_ab1), .a2b2(din_9_ab2),
  .a3b0(din_10_ab0), .a3b1(din_10_ab1), .a3b2(din_10_ab2),
  .a4b0(din_11_ab0), .a4b1(din_11_ab1),
  .a5b0(din_12_ab0), .a5b1(din_12_ab1),
  .a6b0(din_13_ab0),
  .a7b0(din_14_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_8_calc (
  .clk(clk), .p(addr_1_8),
  .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
  .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2), .a1b3(din_9_ab3),
  .a2b0(din_10_ab0), .a2b1(din_10_ab1), .a2b2(din_10_ab2),
  .a3b0(din_11_ab0), .a3b1(din_11_ab1), .a3b2(din_11_ab2),
  .a4b0(din_12_ab0), .a4b1(din_12_ab1),
  .a5b0(din_13_ab0), .a5b1(din_13_ab1),
  .a6b0(din_14_ab0),
  .a7b0(din_15_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_9_calc (
  .clk(clk), .p(addr_1_9),
  .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
  .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2), .a1b3(din_10_ab3),
  .a2b0(din_11_ab0), .a2b1(din_11_ab1), .a2b2(din_11_ab2),
  .a3b0(din_12_ab0), .a3b1(din_12_ab1), .a3b2(din_12_ab2),
  .a4b0(din_13_ab0), .a4b1(din_13_ab1),
  .a5b0(din_14_ab0), .a5b1(din_14_ab1),
  .a6b0(din_15_ab0),
  .a7b0(din_16_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_10_calc (
  .clk(clk), .p(addr_1_10),
  .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
  .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2), .a1b3(din_11_ab3),
  .a2b0(din_12_ab0), .a2b1(din_12_ab1), .a2b2(din_12_ab2),
  .a3b0(din_13_ab0), .a3b1(din_13_ab1), .a3b2(din_13_ab2),
  .a4b0(din_14_ab0), .a4b1(din_14_ab1),
  .a5b0(din_15_ab0), .a5b1(din_15_ab1),
  .a6b0(din_16_ab0),
  .a7b0(din_17_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_11_calc (
  .clk(clk), .p(addr_1_11),
  .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
  .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2), .a1b3(din_12_ab3),
  .a2b0(din_13_ab0), .a2b1(din_13_ab1), .a2b2(din_13_ab2),
  .a3b0(din_14_ab0), .a3b1(din_14_ab1), .a3b2(din_14_ab2),
  .a4b0(din_15_ab0), .a4b1(din_15_ab1),
  .a5b0(din_16_ab0), .a5b1(din_16_ab1),
  .a6b0(din_17_ab0),
  .a7b0(din_18_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_12_calc (
  .clk(clk), .p(addr_1_12),
  .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
  .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2), .a1b3(din_13_ab3),
  .a2b0(din_14_ab0), .a2b1(din_14_ab1), .a2b2(din_14_ab2),
  .a3b0(din_15_ab0), .a3b1(din_15_ab1), .a3b2(din_15_ab2),
  .a4b0(din_16_ab0), .a4b1(din_16_ab1),
  .a5b0(din_17_ab0), .a5b1(din_17_ab1),
  .a6b0(din_18_ab0),
  .a7b0(din_19_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_13_calc (
  .clk(clk), .p(addr_1_13),
  .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
  .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2), .a1b3(din_14_ab3),
  .a2b0(din_15_ab0), .a2b1(din_15_ab1), .a2b2(din_15_ab2),
  .a3b0(din_16_ab0), .a3b1(din_16_ab1), .a3b2(din_16_ab2),
  .a4b0(din_17_ab0), .a4b1(din_17_ab1),
  .a5b0(din_18_ab0), .a5b1(din_18_ab1),
  .a6b0(din_19_ab0),
  .a7b0(din_20_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_14_calc (
  .clk(clk), .p(addr_1_14),
  .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
  .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2), .a1b3(din_15_ab3),
  .a2b0(din_16_ab0), .a2b1(din_16_ab1), .a2b2(din_16_ab2),
  .a3b0(din_17_ab0), .a3b1(din_17_ab1), .a3b2(din_17_ab2),
  .a4b0(din_18_ab0), .a4b1(din_18_ab1),
  .a5b0(din_19_ab0), .a5b1(din_19_ab1),
  .a6b0(din_20_ab0),
  .a7b0(din_21_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(13)
) addr_1_15_calc (
  .clk(clk), .p(addr_1_15),
  .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
  .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2), .a1b3(din_16_ab3),
  .a2b0(din_17_ab0), .a2b1(din_17_ab1), .a2b2(din_17_ab2),
  .a3b0(din_18_ab0), .a3b1(din_18_ab1), .a3b2(din_18_ab2),
  .a4b0(din_19_ab0), .a4b1(din_19_ab1),
  .a5b0(din_20_ab0), .a5b1(din_20_ab1),
  .a6b0(din_21_ab0),
  .a7b0(din_22_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_0_calc (
  .clk(clk), .p(addr_2_0),
  .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
  .a1b0(din_1_ab0), .a1b1(din_1_ab1), .a1b2(din_1_ab2), .a1b3(din_1_ab3),
  .a2b0(din_2_ab0), .a2b1(din_2_ab1), .a2b2(din_2_ab2),
  .a3b0(din_3_ab0), .a3b1(din_3_ab1), .a3b2(din_3_ab2),
  .a4b0(din_4_ab0), .a4b1(din_4_ab1),
  .a5b0(din_5_ab0), .a5b1(din_5_ab1),
  .a6b0(din_6_ab0),
  .a7b0(din_7_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_1_calc (
  .clk(clk), .p(addr_2_1),
  .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
  .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2), .a1b3(din_2_ab3),
  .a2b0(din_3_ab0), .a2b1(din_3_ab1), .a2b2(din_3_ab2),
  .a3b0(din_4_ab0), .a3b1(din_4_ab1), .a3b2(din_4_ab2),
  .a4b0(din_5_ab0), .a4b1(din_5_ab1),
  .a5b0(din_6_ab0), .a5b1(din_6_ab1),
  .a6b0(din_7_ab0),
  .a7b0(din_8_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_2_calc (
  .clk(clk), .p(addr_2_2),
  .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
  .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2), .a1b3(din_3_ab3),
  .a2b0(din_4_ab0), .a2b1(din_4_ab1), .a2b2(din_4_ab2),
  .a3b0(din_5_ab0), .a3b1(din_5_ab1), .a3b2(din_5_ab2),
  .a4b0(din_6_ab0), .a4b1(din_6_ab1),
  .a5b0(din_7_ab0), .a5b1(din_7_ab1),
  .a6b0(din_8_ab0),
  .a7b0(din_9_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_3_calc (
  .clk(clk), .p(addr_2_3),
  .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
  .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2), .a1b3(din_4_ab3),
  .a2b0(din_5_ab0), .a2b1(din_5_ab1), .a2b2(din_5_ab2),
  .a3b0(din_6_ab0), .a3b1(din_6_ab1), .a3b2(din_6_ab2),
  .a4b0(din_7_ab0), .a4b1(din_7_ab1),
  .a5b0(din_8_ab0), .a5b1(din_8_ab1),
  .a6b0(din_9_ab0),
  .a7b0(din_10_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_4_calc (
  .clk(clk), .p(addr_2_4),
  .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
  .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2), .a1b3(din_5_ab3),
  .a2b0(din_6_ab0), .a2b1(din_6_ab1), .a2b2(din_6_ab2),
  .a3b0(din_7_ab0), .a3b1(din_7_ab1), .a3b2(din_7_ab2),
  .a4b0(din_8_ab0), .a4b1(din_8_ab1),
  .a5b0(din_9_ab0), .a5b1(din_9_ab1),
  .a6b0(din_10_ab0),
  .a7b0(din_11_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_5_calc (
  .clk(clk), .p(addr_2_5),
  .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
  .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2), .a1b3(din_6_ab3),
  .a2b0(din_7_ab0), .a2b1(din_7_ab1), .a2b2(din_7_ab2),
  .a3b0(din_8_ab0), .a3b1(din_8_ab1), .a3b2(din_8_ab2),
  .a4b0(din_9_ab0), .a4b1(din_9_ab1),
  .a5b0(din_10_ab0), .a5b1(din_10_ab1),
  .a6b0(din_11_ab0),
  .a7b0(din_12_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_6_calc (
  .clk(clk), .p(addr_2_6),
  .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
  .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2), .a1b3(din_7_ab3),
  .a2b0(din_8_ab0), .a2b1(din_8_ab1), .a2b2(din_8_ab2),
  .a3b0(din_9_ab0), .a3b1(din_9_ab1), .a3b2(din_9_ab2),
  .a4b0(din_10_ab0), .a4b1(din_10_ab1),
  .a5b0(din_11_ab0), .a5b1(din_11_ab1),
  .a6b0(din_12_ab0),
  .a7b0(din_13_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_7_calc (
  .clk(clk), .p(addr_2_7),
  .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
  .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2), .a1b3(din_8_ab3),
  .a2b0(din_9_ab0), .a2b1(din_9_ab1), .a2b2(din_9_ab2),
  .a3b0(din_10_ab0), .a3b1(din_10_ab1), .a3b2(din_10_ab2),
  .a4b0(din_11_ab0), .a4b1(din_11_ab1),
  .a5b0(din_12_ab0), .a5b1(din_12_ab1),
  .a6b0(din_13_ab0),
  .a7b0(din_14_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_8_calc (
  .clk(clk), .p(addr_2_8),
  .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
  .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2), .a1b3(din_9_ab3),
  .a2b0(din_10_ab0), .a2b1(din_10_ab1), .a2b2(din_10_ab2),
  .a3b0(din_11_ab0), .a3b1(din_11_ab1), .a3b2(din_11_ab2),
  .a4b0(din_12_ab0), .a4b1(din_12_ab1),
  .a5b0(din_13_ab0), .a5b1(din_13_ab1),
  .a6b0(din_14_ab0),
  .a7b0(din_15_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_9_calc (
  .clk(clk), .p(addr_2_9),
  .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
  .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2), .a1b3(din_10_ab3),
  .a2b0(din_11_ab0), .a2b1(din_11_ab1), .a2b2(din_11_ab2),
  .a3b0(din_12_ab0), .a3b1(din_12_ab1), .a3b2(din_12_ab2),
  .a4b0(din_13_ab0), .a4b1(din_13_ab1),
  .a5b0(din_14_ab0), .a5b1(din_14_ab1),
  .a6b0(din_15_ab0),
  .a7b0(din_16_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_10_calc (
  .clk(clk), .p(addr_2_10),
  .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
  .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2), .a1b3(din_11_ab3),
  .a2b0(din_12_ab0), .a2b1(din_12_ab1), .a2b2(din_12_ab2),
  .a3b0(din_13_ab0), .a3b1(din_13_ab1), .a3b2(din_13_ab2),
  .a4b0(din_14_ab0), .a4b1(din_14_ab1),
  .a5b0(din_15_ab0), .a5b1(din_15_ab1),
  .a6b0(din_16_ab0),
  .a7b0(din_17_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_11_calc (
  .clk(clk), .p(addr_2_11),
  .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
  .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2), .a1b3(din_12_ab3),
  .a2b0(din_13_ab0), .a2b1(din_13_ab1), .a2b2(din_13_ab2),
  .a3b0(din_14_ab0), .a3b1(din_14_ab1), .a3b2(din_14_ab2),
  .a4b0(din_15_ab0), .a4b1(din_15_ab1),
  .a5b0(din_16_ab0), .a5b1(din_16_ab1),
  .a6b0(din_17_ab0),
  .a7b0(din_18_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_12_calc (
  .clk(clk), .p(addr_2_12),
  .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
  .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2), .a1b3(din_13_ab3),
  .a2b0(din_14_ab0), .a2b1(din_14_ab1), .a2b2(din_14_ab2),
  .a3b0(din_15_ab0), .a3b1(din_15_ab1), .a3b2(din_15_ab2),
  .a4b0(din_16_ab0), .a4b1(din_16_ab1),
  .a5b0(din_17_ab0), .a5b1(din_17_ab1),
  .a6b0(din_18_ab0),
  .a7b0(din_19_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_13_calc (
  .clk(clk), .p(addr_2_13),
  .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
  .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2), .a1b3(din_14_ab3),
  .a2b0(din_15_ab0), .a2b1(din_15_ab1), .a2b2(din_15_ab2),
  .a3b0(din_16_ab0), .a3b1(din_16_ab1), .a3b2(din_16_ab2),
  .a4b0(din_17_ab0), .a4b1(din_17_ab1),
  .a5b0(din_18_ab0), .a5b1(din_18_ab1),
  .a6b0(din_19_ab0),
  .a7b0(din_20_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_14_calc (
  .clk(clk), .p(addr_2_14),
  .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
  .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2), .a1b3(din_15_ab3),
  .a2b0(din_16_ab0), .a2b1(din_16_ab1), .a2b2(din_16_ab2),
  .a3b0(din_17_ab0), .a3b1(din_17_ab1), .a3b2(din_17_ab2),
  .a4b0(din_18_ab0), .a4b1(din_18_ab1),
  .a5b0(din_19_ab0), .a5b1(din_19_ab1),
  .a6b0(din_20_ab0),
  .a7b0(din_21_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(13)
) addr_2_15_calc (
  .clk(clk), .p(addr_2_15),
  .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
  .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2), .a1b3(din_16_ab3),
  .a2b0(din_17_ab0), .a2b1(din_17_ab1), .a2b2(din_17_ab2),
  .a3b0(din_18_ab0), .a3b1(din_18_ab1), .a3b2(din_18_ab2),
  .a4b0(din_19_ab0), .a4b1(din_19_ab1),
  .a5b0(din_20_ab0), .a5b1(din_20_ab1),
  .a6b0(din_21_ab0),
  .a7b0(din_22_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_0_calc (
  .clk(clk), .p(addr_3_0),
  .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
  .a1b0(din_1_ab0), .a1b1(din_1_ab1), .a1b2(din_1_ab2), .a1b3(din_1_ab3),
  .a2b0(din_2_ab0), .a2b1(din_2_ab1), .a2b2(din_2_ab2),
  .a3b0(din_3_ab0), .a3b1(din_3_ab1), .a3b2(din_3_ab2),
  .a4b0(din_4_ab0), .a4b1(din_4_ab1),
  .a5b0(din_5_ab0), .a5b1(din_5_ab1),
  .a6b0(din_6_ab0),
  .a7b0(din_7_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_1_calc (
  .clk(clk), .p(addr_3_1),
  .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
  .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2), .a1b3(din_2_ab3),
  .a2b0(din_3_ab0), .a2b1(din_3_ab1), .a2b2(din_3_ab2),
  .a3b0(din_4_ab0), .a3b1(din_4_ab1), .a3b2(din_4_ab2),
  .a4b0(din_5_ab0), .a4b1(din_5_ab1),
  .a5b0(din_6_ab0), .a5b1(din_6_ab1),
  .a6b0(din_7_ab0),
  .a7b0(din_8_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_2_calc (
  .clk(clk), .p(addr_3_2),
  .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
  .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2), .a1b3(din_3_ab3),
  .a2b0(din_4_ab0), .a2b1(din_4_ab1), .a2b2(din_4_ab2),
  .a3b0(din_5_ab0), .a3b1(din_5_ab1), .a3b2(din_5_ab2),
  .a4b0(din_6_ab0), .a4b1(din_6_ab1),
  .a5b0(din_7_ab0), .a5b1(din_7_ab1),
  .a6b0(din_8_ab0),
  .a7b0(din_9_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_3_calc (
  .clk(clk), .p(addr_3_3),
  .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
  .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2), .a1b3(din_4_ab3),
  .a2b0(din_5_ab0), .a2b1(din_5_ab1), .a2b2(din_5_ab2),
  .a3b0(din_6_ab0), .a3b1(din_6_ab1), .a3b2(din_6_ab2),
  .a4b0(din_7_ab0), .a4b1(din_7_ab1),
  .a5b0(din_8_ab0), .a5b1(din_8_ab1),
  .a6b0(din_9_ab0),
  .a7b0(din_10_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_4_calc (
  .clk(clk), .p(addr_3_4),
  .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
  .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2), .a1b3(din_5_ab3),
  .a2b0(din_6_ab0), .a2b1(din_6_ab1), .a2b2(din_6_ab2),
  .a3b0(din_7_ab0), .a3b1(din_7_ab1), .a3b2(din_7_ab2),
  .a4b0(din_8_ab0), .a4b1(din_8_ab1),
  .a5b0(din_9_ab0), .a5b1(din_9_ab1),
  .a6b0(din_10_ab0),
  .a7b0(din_11_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_5_calc (
  .clk(clk), .p(addr_3_5),
  .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
  .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2), .a1b3(din_6_ab3),
  .a2b0(din_7_ab0), .a2b1(din_7_ab1), .a2b2(din_7_ab2),
  .a3b0(din_8_ab0), .a3b1(din_8_ab1), .a3b2(din_8_ab2),
  .a4b0(din_9_ab0), .a4b1(din_9_ab1),
  .a5b0(din_10_ab0), .a5b1(din_10_ab1),
  .a6b0(din_11_ab0),
  .a7b0(din_12_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_6_calc (
  .clk(clk), .p(addr_3_6),
  .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
  .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2), .a1b3(din_7_ab3),
  .a2b0(din_8_ab0), .a2b1(din_8_ab1), .a2b2(din_8_ab2),
  .a3b0(din_9_ab0), .a3b1(din_9_ab1), .a3b2(din_9_ab2),
  .a4b0(din_10_ab0), .a4b1(din_10_ab1),
  .a5b0(din_11_ab0), .a5b1(din_11_ab1),
  .a6b0(din_12_ab0),
  .a7b0(din_13_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_7_calc (
  .clk(clk), .p(addr_3_7),
  .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
  .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2), .a1b3(din_8_ab3),
  .a2b0(din_9_ab0), .a2b1(din_9_ab1), .a2b2(din_9_ab2),
  .a3b0(din_10_ab0), .a3b1(din_10_ab1), .a3b2(din_10_ab2),
  .a4b0(din_11_ab0), .a4b1(din_11_ab1),
  .a5b0(din_12_ab0), .a5b1(din_12_ab1),
  .a6b0(din_13_ab0),
  .a7b0(din_14_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_8_calc (
  .clk(clk), .p(addr_3_8),
  .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
  .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2), .a1b3(din_9_ab3),
  .a2b0(din_10_ab0), .a2b1(din_10_ab1), .a2b2(din_10_ab2),
  .a3b0(din_11_ab0), .a3b1(din_11_ab1), .a3b2(din_11_ab2),
  .a4b0(din_12_ab0), .a4b1(din_12_ab1),
  .a5b0(din_13_ab0), .a5b1(din_13_ab1),
  .a6b0(din_14_ab0),
  .a7b0(din_15_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_9_calc (
  .clk(clk), .p(addr_3_9),
  .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
  .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2), .a1b3(din_10_ab3),
  .a2b0(din_11_ab0), .a2b1(din_11_ab1), .a2b2(din_11_ab2),
  .a3b0(din_12_ab0), .a3b1(din_12_ab1), .a3b2(din_12_ab2),
  .a4b0(din_13_ab0), .a4b1(din_13_ab1),
  .a5b0(din_14_ab0), .a5b1(din_14_ab1),
  .a6b0(din_15_ab0),
  .a7b0(din_16_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_10_calc (
  .clk(clk), .p(addr_3_10),
  .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
  .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2), .a1b3(din_11_ab3),
  .a2b0(din_12_ab0), .a2b1(din_12_ab1), .a2b2(din_12_ab2),
  .a3b0(din_13_ab0), .a3b1(din_13_ab1), .a3b2(din_13_ab2),
  .a4b0(din_14_ab0), .a4b1(din_14_ab1),
  .a5b0(din_15_ab0), .a5b1(din_15_ab1),
  .a6b0(din_16_ab0),
  .a7b0(din_17_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_11_calc (
  .clk(clk), .p(addr_3_11),
  .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
  .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2), .a1b3(din_12_ab3),
  .a2b0(din_13_ab0), .a2b1(din_13_ab1), .a2b2(din_13_ab2),
  .a3b0(din_14_ab0), .a3b1(din_14_ab1), .a3b2(din_14_ab2),
  .a4b0(din_15_ab0), .a4b1(din_15_ab1),
  .a5b0(din_16_ab0), .a5b1(din_16_ab1),
  .a6b0(din_17_ab0),
  .a7b0(din_18_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_12_calc (
  .clk(clk), .p(addr_3_12),
  .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
  .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2), .a1b3(din_13_ab3),
  .a2b0(din_14_ab0), .a2b1(din_14_ab1), .a2b2(din_14_ab2),
  .a3b0(din_15_ab0), .a3b1(din_15_ab1), .a3b2(din_15_ab2),
  .a4b0(din_16_ab0), .a4b1(din_16_ab1),
  .a5b0(din_17_ab0), .a5b1(din_17_ab1),
  .a6b0(din_18_ab0),
  .a7b0(din_19_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_13_calc (
  .clk(clk), .p(addr_3_13),
  .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
  .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2), .a1b3(din_14_ab3),
  .a2b0(din_15_ab0), .a2b1(din_15_ab1), .a2b2(din_15_ab2),
  .a3b0(din_16_ab0), .a3b1(din_16_ab1), .a3b2(din_16_ab2),
  .a4b0(din_17_ab0), .a4b1(din_17_ab1),
  .a5b0(din_18_ab0), .a5b1(din_18_ab1),
  .a6b0(din_19_ab0),
  .a7b0(din_20_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_14_calc (
  .clk(clk), .p(addr_3_14),
  .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
  .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2), .a1b3(din_15_ab3),
  .a2b0(din_16_ab0), .a2b1(din_16_ab1), .a2b2(din_16_ab2),
  .a3b0(din_17_ab0), .a3b1(din_17_ab1), .a3b2(din_17_ab2),
  .a4b0(din_18_ab0), .a4b1(din_18_ab1),
  .a5b0(din_19_ab0), .a5b1(din_19_ab1),
  .a6b0(din_20_ab0),
  .a7b0(din_21_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffffff000000),
	.NBITS(13)
) addr_3_15_calc (
  .clk(clk), .p(addr_3_15),
  .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
  .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2), .a1b3(din_16_ab3),
  .a2b0(din_17_ab0), .a2b1(din_17_ab1), .a2b2(din_17_ab2),
  .a3b0(din_18_ab0), .a3b1(din_18_ab1), .a3b2(din_18_ab2),
  .a4b0(din_19_ab0), .a4b1(din_19_ab1),
  .a5b0(din_20_ab0), .a5b1(din_20_ab1),
  .a6b0(din_21_ab0),
  .a7b0(din_22_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_0_calc (
  .clk(clk), .p(addr_4_0),
  .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
  .a1b0(din_1_ab0), .a1b1(din_1_ab1), .a1b2(din_1_ab2), .a1b3(din_1_ab3),
  .a2b0(din_2_ab0), .a2b1(din_2_ab1), .a2b2(din_2_ab2),
  .a3b0(din_3_ab0), .a3b1(din_3_ab1), .a3b2(din_3_ab2),
  .a4b0(din_4_ab0), .a4b1(din_4_ab1),
  .a5b0(din_5_ab0), .a5b1(din_5_ab1),
  .a6b0(din_6_ab0),
  .a7b0(din_7_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_1_calc (
  .clk(clk), .p(addr_4_1),
  .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
  .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2), .a1b3(din_2_ab3),
  .a2b0(din_3_ab0), .a2b1(din_3_ab1), .a2b2(din_3_ab2),
  .a3b0(din_4_ab0), .a3b1(din_4_ab1), .a3b2(din_4_ab2),
  .a4b0(din_5_ab0), .a4b1(din_5_ab1),
  .a5b0(din_6_ab0), .a5b1(din_6_ab1),
  .a6b0(din_7_ab0),
  .a7b0(din_8_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_2_calc (
  .clk(clk), .p(addr_4_2),
  .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
  .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2), .a1b3(din_3_ab3),
  .a2b0(din_4_ab0), .a2b1(din_4_ab1), .a2b2(din_4_ab2),
  .a3b0(din_5_ab0), .a3b1(din_5_ab1), .a3b2(din_5_ab2),
  .a4b0(din_6_ab0), .a4b1(din_6_ab1),
  .a5b0(din_7_ab0), .a5b1(din_7_ab1),
  .a6b0(din_8_ab0),
  .a7b0(din_9_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_3_calc (
  .clk(clk), .p(addr_4_3),
  .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
  .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2), .a1b3(din_4_ab3),
  .a2b0(din_5_ab0), .a2b1(din_5_ab1), .a2b2(din_5_ab2),
  .a3b0(din_6_ab0), .a3b1(din_6_ab1), .a3b2(din_6_ab2),
  .a4b0(din_7_ab0), .a4b1(din_7_ab1),
  .a5b0(din_8_ab0), .a5b1(din_8_ab1),
  .a6b0(din_9_ab0),
  .a7b0(din_10_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_4_calc (
  .clk(clk), .p(addr_4_4),
  .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
  .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2), .a1b3(din_5_ab3),
  .a2b0(din_6_ab0), .a2b1(din_6_ab1), .a2b2(din_6_ab2),
  .a3b0(din_7_ab0), .a3b1(din_7_ab1), .a3b2(din_7_ab2),
  .a4b0(din_8_ab0), .a4b1(din_8_ab1),
  .a5b0(din_9_ab0), .a5b1(din_9_ab1),
  .a6b0(din_10_ab0),
  .a7b0(din_11_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_5_calc (
  .clk(clk), .p(addr_4_5),
  .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
  .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2), .a1b3(din_6_ab3),
  .a2b0(din_7_ab0), .a2b1(din_7_ab1), .a2b2(din_7_ab2),
  .a3b0(din_8_ab0), .a3b1(din_8_ab1), .a3b2(din_8_ab2),
  .a4b0(din_9_ab0), .a4b1(din_9_ab1),
  .a5b0(din_10_ab0), .a5b1(din_10_ab1),
  .a6b0(din_11_ab0),
  .a7b0(din_12_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_6_calc (
  .clk(clk), .p(addr_4_6),
  .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
  .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2), .a1b3(din_7_ab3),
  .a2b0(din_8_ab0), .a2b1(din_8_ab1), .a2b2(din_8_ab2),
  .a3b0(din_9_ab0), .a3b1(din_9_ab1), .a3b2(din_9_ab2),
  .a4b0(din_10_ab0), .a4b1(din_10_ab1),
  .a5b0(din_11_ab0), .a5b1(din_11_ab1),
  .a6b0(din_12_ab0),
  .a7b0(din_13_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_7_calc (
  .clk(clk), .p(addr_4_7),
  .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
  .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2), .a1b3(din_8_ab3),
  .a2b0(din_9_ab0), .a2b1(din_9_ab1), .a2b2(din_9_ab2),
  .a3b0(din_10_ab0), .a3b1(din_10_ab1), .a3b2(din_10_ab2),
  .a4b0(din_11_ab0), .a4b1(din_11_ab1),
  .a5b0(din_12_ab0), .a5b1(din_12_ab1),
  .a6b0(din_13_ab0),
  .a7b0(din_14_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_8_calc (
  .clk(clk), .p(addr_4_8),
  .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
  .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2), .a1b3(din_9_ab3),
  .a2b0(din_10_ab0), .a2b1(din_10_ab1), .a2b2(din_10_ab2),
  .a3b0(din_11_ab0), .a3b1(din_11_ab1), .a3b2(din_11_ab2),
  .a4b0(din_12_ab0), .a4b1(din_12_ab1),
  .a5b0(din_13_ab0), .a5b1(din_13_ab1),
  .a6b0(din_14_ab0),
  .a7b0(din_15_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_9_calc (
  .clk(clk), .p(addr_4_9),
  .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
  .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2), .a1b3(din_10_ab3),
  .a2b0(din_11_ab0), .a2b1(din_11_ab1), .a2b2(din_11_ab2),
  .a3b0(din_12_ab0), .a3b1(din_12_ab1), .a3b2(din_12_ab2),
  .a4b0(din_13_ab0), .a4b1(din_13_ab1),
  .a5b0(din_14_ab0), .a5b1(din_14_ab1),
  .a6b0(din_15_ab0),
  .a7b0(din_16_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_10_calc (
  .clk(clk), .p(addr_4_10),
  .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
  .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2), .a1b3(din_11_ab3),
  .a2b0(din_12_ab0), .a2b1(din_12_ab1), .a2b2(din_12_ab2),
  .a3b0(din_13_ab0), .a3b1(din_13_ab1), .a3b2(din_13_ab2),
  .a4b0(din_14_ab0), .a4b1(din_14_ab1),
  .a5b0(din_15_ab0), .a5b1(din_15_ab1),
  .a6b0(din_16_ab0),
  .a7b0(din_17_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_11_calc (
  .clk(clk), .p(addr_4_11),
  .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
  .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2), .a1b3(din_12_ab3),
  .a2b0(din_13_ab0), .a2b1(din_13_ab1), .a2b2(din_13_ab2),
  .a3b0(din_14_ab0), .a3b1(din_14_ab1), .a3b2(din_14_ab2),
  .a4b0(din_15_ab0), .a4b1(din_15_ab1),
  .a5b0(din_16_ab0), .a5b1(din_16_ab1),
  .a6b0(din_17_ab0),
  .a7b0(din_18_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_12_calc (
  .clk(clk), .p(addr_4_12),
  .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
  .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2), .a1b3(din_13_ab3),
  .a2b0(din_14_ab0), .a2b1(din_14_ab1), .a2b2(din_14_ab2),
  .a3b0(din_15_ab0), .a3b1(din_15_ab1), .a3b2(din_15_ab2),
  .a4b0(din_16_ab0), .a4b1(din_16_ab1),
  .a5b0(din_17_ab0), .a5b1(din_17_ab1),
  .a6b0(din_18_ab0),
  .a7b0(din_19_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_13_calc (
  .clk(clk), .p(addr_4_13),
  .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
  .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2), .a1b3(din_14_ab3),
  .a2b0(din_15_ab0), .a2b1(din_15_ab1), .a2b2(din_15_ab2),
  .a3b0(din_16_ab0), .a3b1(din_16_ab1), .a3b2(din_16_ab2),
  .a4b0(din_17_ab0), .a4b1(din_17_ab1),
  .a5b0(din_18_ab0), .a5b1(din_18_ab1),
  .a6b0(din_19_ab0),
  .a7b0(din_20_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_14_calc (
  .clk(clk), .p(addr_4_14),
  .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
  .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2), .a1b3(din_15_ab3),
  .a2b0(din_16_ab0), .a2b1(din_16_ab1), .a2b2(din_16_ab2),
  .a3b0(din_17_ab0), .a3b1(din_17_ab1), .a3b2(din_17_ab2),
  .a4b0(din_18_ab0), .a4b1(din_18_ab1),
  .a5b0(din_19_ab0), .a5b1(din_19_ab1),
  .a6b0(din_20_ab0),
  .a7b0(din_21_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffffff00000000),
	.NBITS(13)
) addr_4_15_calc (
  .clk(clk), .p(addr_4_15),
  .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
  .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2), .a1b3(din_16_ab3),
  .a2b0(din_17_ab0), .a2b1(din_17_ab1), .a2b2(din_17_ab2),
  .a3b0(din_18_ab0), .a3b1(din_18_ab1), .a3b2(din_18_ab2),
  .a4b0(din_19_ab0), .a4b1(din_19_ab1),
  .a5b0(din_20_ab0), .a5b1(din_20_ab1),
  .a6b0(din_21_ab0),
  .a7b0(din_22_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_0_calc (
  .clk(clk), .p(addr_5_0),
  .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
  .a1b0(din_1_ab0), .a1b1(din_1_ab1), .a1b2(din_1_ab2), .a1b3(din_1_ab3),
  .a2b0(din_2_ab0), .a2b1(din_2_ab1), .a2b2(din_2_ab2),
  .a3b0(din_3_ab0), .a3b1(din_3_ab1), .a3b2(din_3_ab2),
  .a4b0(din_4_ab0), .a4b1(din_4_ab1),
  .a5b0(din_5_ab0), .a5b1(din_5_ab1),
  .a6b0(din_6_ab0),
  .a7b0(din_7_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_1_calc (
  .clk(clk), .p(addr_5_1),
  .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
  .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2), .a1b3(din_2_ab3),
  .a2b0(din_3_ab0), .a2b1(din_3_ab1), .a2b2(din_3_ab2),
  .a3b0(din_4_ab0), .a3b1(din_4_ab1), .a3b2(din_4_ab2),
  .a4b0(din_5_ab0), .a4b1(din_5_ab1),
  .a5b0(din_6_ab0), .a5b1(din_6_ab1),
  .a6b0(din_7_ab0),
  .a7b0(din_8_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_2_calc (
  .clk(clk), .p(addr_5_2),
  .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
  .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2), .a1b3(din_3_ab3),
  .a2b0(din_4_ab0), .a2b1(din_4_ab1), .a2b2(din_4_ab2),
  .a3b0(din_5_ab0), .a3b1(din_5_ab1), .a3b2(din_5_ab2),
  .a4b0(din_6_ab0), .a4b1(din_6_ab1),
  .a5b0(din_7_ab0), .a5b1(din_7_ab1),
  .a6b0(din_8_ab0),
  .a7b0(din_9_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_3_calc (
  .clk(clk), .p(addr_5_3),
  .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
  .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2), .a1b3(din_4_ab3),
  .a2b0(din_5_ab0), .a2b1(din_5_ab1), .a2b2(din_5_ab2),
  .a3b0(din_6_ab0), .a3b1(din_6_ab1), .a3b2(din_6_ab2),
  .a4b0(din_7_ab0), .a4b1(din_7_ab1),
  .a5b0(din_8_ab0), .a5b1(din_8_ab1),
  .a6b0(din_9_ab0),
  .a7b0(din_10_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_4_calc (
  .clk(clk), .p(addr_5_4),
  .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
  .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2), .a1b3(din_5_ab3),
  .a2b0(din_6_ab0), .a2b1(din_6_ab1), .a2b2(din_6_ab2),
  .a3b0(din_7_ab0), .a3b1(din_7_ab1), .a3b2(din_7_ab2),
  .a4b0(din_8_ab0), .a4b1(din_8_ab1),
  .a5b0(din_9_ab0), .a5b1(din_9_ab1),
  .a6b0(din_10_ab0),
  .a7b0(din_11_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_5_calc (
  .clk(clk), .p(addr_5_5),
  .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
  .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2), .a1b3(din_6_ab3),
  .a2b0(din_7_ab0), .a2b1(din_7_ab1), .a2b2(din_7_ab2),
  .a3b0(din_8_ab0), .a3b1(din_8_ab1), .a3b2(din_8_ab2),
  .a4b0(din_9_ab0), .a4b1(din_9_ab1),
  .a5b0(din_10_ab0), .a5b1(din_10_ab1),
  .a6b0(din_11_ab0),
  .a7b0(din_12_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_6_calc (
  .clk(clk), .p(addr_5_6),
  .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
  .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2), .a1b3(din_7_ab3),
  .a2b0(din_8_ab0), .a2b1(din_8_ab1), .a2b2(din_8_ab2),
  .a3b0(din_9_ab0), .a3b1(din_9_ab1), .a3b2(din_9_ab2),
  .a4b0(din_10_ab0), .a4b1(din_10_ab1),
  .a5b0(din_11_ab0), .a5b1(din_11_ab1),
  .a6b0(din_12_ab0),
  .a7b0(din_13_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_7_calc (
  .clk(clk), .p(addr_5_7),
  .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
  .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2), .a1b3(din_8_ab3),
  .a2b0(din_9_ab0), .a2b1(din_9_ab1), .a2b2(din_9_ab2),
  .a3b0(din_10_ab0), .a3b1(din_10_ab1), .a3b2(din_10_ab2),
  .a4b0(din_11_ab0), .a4b1(din_11_ab1),
  .a5b0(din_12_ab0), .a5b1(din_12_ab1),
  .a6b0(din_13_ab0),
  .a7b0(din_14_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_8_calc (
  .clk(clk), .p(addr_5_8),
  .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
  .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2), .a1b3(din_9_ab3),
  .a2b0(din_10_ab0), .a2b1(din_10_ab1), .a2b2(din_10_ab2),
  .a3b0(din_11_ab0), .a3b1(din_11_ab1), .a3b2(din_11_ab2),
  .a4b0(din_12_ab0), .a4b1(din_12_ab1),
  .a5b0(din_13_ab0), .a5b1(din_13_ab1),
  .a6b0(din_14_ab0),
  .a7b0(din_15_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_9_calc (
  .clk(clk), .p(addr_5_9),
  .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
  .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2), .a1b3(din_10_ab3),
  .a2b0(din_11_ab0), .a2b1(din_11_ab1), .a2b2(din_11_ab2),
  .a3b0(din_12_ab0), .a3b1(din_12_ab1), .a3b2(din_12_ab2),
  .a4b0(din_13_ab0), .a4b1(din_13_ab1),
  .a5b0(din_14_ab0), .a5b1(din_14_ab1),
  .a6b0(din_15_ab0),
  .a7b0(din_16_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_10_calc (
  .clk(clk), .p(addr_5_10),
  .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
  .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2), .a1b3(din_11_ab3),
  .a2b0(din_12_ab0), .a2b1(din_12_ab1), .a2b2(din_12_ab2),
  .a3b0(din_13_ab0), .a3b1(din_13_ab1), .a3b2(din_13_ab2),
  .a4b0(din_14_ab0), .a4b1(din_14_ab1),
  .a5b0(din_15_ab0), .a5b1(din_15_ab1),
  .a6b0(din_16_ab0),
  .a7b0(din_17_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_11_calc (
  .clk(clk), .p(addr_5_11),
  .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
  .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2), .a1b3(din_12_ab3),
  .a2b0(din_13_ab0), .a2b1(din_13_ab1), .a2b2(din_13_ab2),
  .a3b0(din_14_ab0), .a3b1(din_14_ab1), .a3b2(din_14_ab2),
  .a4b0(din_15_ab0), .a4b1(din_15_ab1),
  .a5b0(din_16_ab0), .a5b1(din_16_ab1),
  .a6b0(din_17_ab0),
  .a7b0(din_18_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_12_calc (
  .clk(clk), .p(addr_5_12),
  .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
  .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2), .a1b3(din_13_ab3),
  .a2b0(din_14_ab0), .a2b1(din_14_ab1), .a2b2(din_14_ab2),
  .a3b0(din_15_ab0), .a3b1(din_15_ab1), .a3b2(din_15_ab2),
  .a4b0(din_16_ab0), .a4b1(din_16_ab1),
  .a5b0(din_17_ab0), .a5b1(din_17_ab1),
  .a6b0(din_18_ab0),
  .a7b0(din_19_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_13_calc (
  .clk(clk), .p(addr_5_13),
  .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
  .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2), .a1b3(din_14_ab3),
  .a2b0(din_15_ab0), .a2b1(din_15_ab1), .a2b2(din_15_ab2),
  .a3b0(din_16_ab0), .a3b1(din_16_ab1), .a3b2(din_16_ab2),
  .a4b0(din_17_ab0), .a4b1(din_17_ab1),
  .a5b0(din_18_ab0), .a5b1(din_18_ab1),
  .a6b0(din_19_ab0),
  .a7b0(din_20_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_14_calc (
  .clk(clk), .p(addr_5_14),
  .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
  .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2), .a1b3(din_15_ab3),
  .a2b0(din_16_ab0), .a2b1(din_16_ab1), .a2b2(din_16_ab2),
  .a3b0(din_17_ab0), .a3b1(din_17_ab1), .a3b2(din_17_ab2),
  .a4b0(din_18_ab0), .a4b1(din_18_ab1),
  .a5b0(din_19_ab0), .a5b1(din_19_ab1),
  .a6b0(din_20_ab0),
  .a7b0(din_21_ab0)
);

acc_hash # (
	.ANDMSK(64'hffffff0000000000),
	.NBITS(12)
) addr_5_15_calc (
  .clk(clk), .p(addr_5_15),
  .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
  .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2), .a1b3(din_16_ab3),
  .a2b0(din_17_ab0), .a2b1(din_17_ab1), .a2b2(din_17_ab2),
  .a3b0(din_18_ab0), .a3b1(din_18_ab1), .a3b2(din_18_ab2),
  .a4b0(din_19_ab0), .a4b1(din_19_ab1),
  .a5b0(din_20_ab0), .a5b1(din_20_ab1),
  .a6b0(din_21_ab0),
  .a7b0(din_22_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_0_calc (
  .clk(clk), .p(addr_6_0),
  .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
  .a1b0(din_1_ab0), .a1b1(din_1_ab1), .a1b2(din_1_ab2), .a1b3(din_1_ab3),
  .a2b0(din_2_ab0), .a2b1(din_2_ab1), .a2b2(din_2_ab2),
  .a3b0(din_3_ab0), .a3b1(din_3_ab1), .a3b2(din_3_ab2),
  .a4b0(din_4_ab0), .a4b1(din_4_ab1),
  .a5b0(din_5_ab0), .a5b1(din_5_ab1),
  .a6b0(din_6_ab0),
  .a7b0(din_7_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_1_calc (
  .clk(clk), .p(addr_6_1),
  .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
  .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2), .a1b3(din_2_ab3),
  .a2b0(din_3_ab0), .a2b1(din_3_ab1), .a2b2(din_3_ab2),
  .a3b0(din_4_ab0), .a3b1(din_4_ab1), .a3b2(din_4_ab2),
  .a4b0(din_5_ab0), .a4b1(din_5_ab1),
  .a5b0(din_6_ab0), .a5b1(din_6_ab1),
  .a6b0(din_7_ab0),
  .a7b0(din_8_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_2_calc (
  .clk(clk), .p(addr_6_2),
  .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
  .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2), .a1b3(din_3_ab3),
  .a2b0(din_4_ab0), .a2b1(din_4_ab1), .a2b2(din_4_ab2),
  .a3b0(din_5_ab0), .a3b1(din_5_ab1), .a3b2(din_5_ab2),
  .a4b0(din_6_ab0), .a4b1(din_6_ab1),
  .a5b0(din_7_ab0), .a5b1(din_7_ab1),
  .a6b0(din_8_ab0),
  .a7b0(din_9_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_3_calc (
  .clk(clk), .p(addr_6_3),
  .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
  .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2), .a1b3(din_4_ab3),
  .a2b0(din_5_ab0), .a2b1(din_5_ab1), .a2b2(din_5_ab2),
  .a3b0(din_6_ab0), .a3b1(din_6_ab1), .a3b2(din_6_ab2),
  .a4b0(din_7_ab0), .a4b1(din_7_ab1),
  .a5b0(din_8_ab0), .a5b1(din_8_ab1),
  .a6b0(din_9_ab0),
  .a7b0(din_10_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_4_calc (
  .clk(clk), .p(addr_6_4),
  .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
  .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2), .a1b3(din_5_ab3),
  .a2b0(din_6_ab0), .a2b1(din_6_ab1), .a2b2(din_6_ab2),
  .a3b0(din_7_ab0), .a3b1(din_7_ab1), .a3b2(din_7_ab2),
  .a4b0(din_8_ab0), .a4b1(din_8_ab1),
  .a5b0(din_9_ab0), .a5b1(din_9_ab1),
  .a6b0(din_10_ab0),
  .a7b0(din_11_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_5_calc (
  .clk(clk), .p(addr_6_5),
  .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
  .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2), .a1b3(din_6_ab3),
  .a2b0(din_7_ab0), .a2b1(din_7_ab1), .a2b2(din_7_ab2),
  .a3b0(din_8_ab0), .a3b1(din_8_ab1), .a3b2(din_8_ab2),
  .a4b0(din_9_ab0), .a4b1(din_9_ab1),
  .a5b0(din_10_ab0), .a5b1(din_10_ab1),
  .a6b0(din_11_ab0),
  .a7b0(din_12_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_6_calc (
  .clk(clk), .p(addr_6_6),
  .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
  .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2), .a1b3(din_7_ab3),
  .a2b0(din_8_ab0), .a2b1(din_8_ab1), .a2b2(din_8_ab2),
  .a3b0(din_9_ab0), .a3b1(din_9_ab1), .a3b2(din_9_ab2),
  .a4b0(din_10_ab0), .a4b1(din_10_ab1),
  .a5b0(din_11_ab0), .a5b1(din_11_ab1),
  .a6b0(din_12_ab0),
  .a7b0(din_13_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_7_calc (
  .clk(clk), .p(addr_6_7),
  .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
  .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2), .a1b3(din_8_ab3),
  .a2b0(din_9_ab0), .a2b1(din_9_ab1), .a2b2(din_9_ab2),
  .a3b0(din_10_ab0), .a3b1(din_10_ab1), .a3b2(din_10_ab2),
  .a4b0(din_11_ab0), .a4b1(din_11_ab1),
  .a5b0(din_12_ab0), .a5b1(din_12_ab1),
  .a6b0(din_13_ab0),
  .a7b0(din_14_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_8_calc (
  .clk(clk), .p(addr_6_8),
  .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
  .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2), .a1b3(din_9_ab3),
  .a2b0(din_10_ab0), .a2b1(din_10_ab1), .a2b2(din_10_ab2),
  .a3b0(din_11_ab0), .a3b1(din_11_ab1), .a3b2(din_11_ab2),
  .a4b0(din_12_ab0), .a4b1(din_12_ab1),
  .a5b0(din_13_ab0), .a5b1(din_13_ab1),
  .a6b0(din_14_ab0),
  .a7b0(din_15_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_9_calc (
  .clk(clk), .p(addr_6_9),
  .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
  .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2), .a1b3(din_10_ab3),
  .a2b0(din_11_ab0), .a2b1(din_11_ab1), .a2b2(din_11_ab2),
  .a3b0(din_12_ab0), .a3b1(din_12_ab1), .a3b2(din_12_ab2),
  .a4b0(din_13_ab0), .a4b1(din_13_ab1),
  .a5b0(din_14_ab0), .a5b1(din_14_ab1),
  .a6b0(din_15_ab0),
  .a7b0(din_16_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_10_calc (
  .clk(clk), .p(addr_6_10),
  .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
  .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2), .a1b3(din_11_ab3),
  .a2b0(din_12_ab0), .a2b1(din_12_ab1), .a2b2(din_12_ab2),
  .a3b0(din_13_ab0), .a3b1(din_13_ab1), .a3b2(din_13_ab2),
  .a4b0(din_14_ab0), .a4b1(din_14_ab1),
  .a5b0(din_15_ab0), .a5b1(din_15_ab1),
  .a6b0(din_16_ab0),
  .a7b0(din_17_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_11_calc (
  .clk(clk), .p(addr_6_11),
  .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
  .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2), .a1b3(din_12_ab3),
  .a2b0(din_13_ab0), .a2b1(din_13_ab1), .a2b2(din_13_ab2),
  .a3b0(din_14_ab0), .a3b1(din_14_ab1), .a3b2(din_14_ab2),
  .a4b0(din_15_ab0), .a4b1(din_15_ab1),
  .a5b0(din_16_ab0), .a5b1(din_16_ab1),
  .a6b0(din_17_ab0),
  .a7b0(din_18_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_12_calc (
  .clk(clk), .p(addr_6_12),
  .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
  .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2), .a1b3(din_13_ab3),
  .a2b0(din_14_ab0), .a2b1(din_14_ab1), .a2b2(din_14_ab2),
  .a3b0(din_15_ab0), .a3b1(din_15_ab1), .a3b2(din_15_ab2),
  .a4b0(din_16_ab0), .a4b1(din_16_ab1),
  .a5b0(din_17_ab0), .a5b1(din_17_ab1),
  .a6b0(din_18_ab0),
  .a7b0(din_19_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_13_calc (
  .clk(clk), .p(addr_6_13),
  .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
  .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2), .a1b3(din_14_ab3),
  .a2b0(din_15_ab0), .a2b1(din_15_ab1), .a2b2(din_15_ab2),
  .a3b0(din_16_ab0), .a3b1(din_16_ab1), .a3b2(din_16_ab2),
  .a4b0(din_17_ab0), .a4b1(din_17_ab1),
  .a5b0(din_18_ab0), .a5b1(din_18_ab1),
  .a6b0(din_19_ab0),
  .a7b0(din_20_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_14_calc (
  .clk(clk), .p(addr_6_14),
  .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
  .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2), .a1b3(din_15_ab3),
  .a2b0(din_16_ab0), .a2b1(din_16_ab1), .a2b2(din_16_ab2),
  .a3b0(din_17_ab0), .a3b1(din_17_ab1), .a3b2(din_17_ab2),
  .a4b0(din_18_ab0), .a4b1(din_18_ab1),
  .a5b0(din_19_ab0), .a5b1(din_19_ab1),
  .a6b0(din_20_ab0),
  .a7b0(din_21_ab0)
);

acc_hash # (
	.ANDMSK(64'hffff000000000000),
	.NBITS(11)
) addr_6_15_calc (
  .clk(clk), .p(addr_6_15),
  .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
  .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2), .a1b3(din_16_ab3),
  .a2b0(din_17_ab0), .a2b1(din_17_ab1), .a2b2(din_17_ab2),
  .a3b0(din_18_ab0), .a3b1(din_18_ab1), .a3b2(din_18_ab2),
  .a4b0(din_19_ab0), .a4b1(din_19_ab1),
  .a5b0(din_20_ab0), .a5b1(din_20_ab1),
  .a6b0(din_21_ab0),
  .a7b0(din_22_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_0_calc (
  .clk(clk), .p(addr_7_0),
  .a0b0(din_0_ab0), .a0b1(din_0_ab1), .a0b2(din_0_ab2), .a0b3(din_0_ab3),
  .a1b0(din_1_ab0), .a1b1(din_1_ab1), .a1b2(din_1_ab2), .a1b3(din_1_ab3),
  .a2b0(din_2_ab0), .a2b1(din_2_ab1), .a2b2(din_2_ab2),
  .a3b0(din_3_ab0), .a3b1(din_3_ab1), .a3b2(din_3_ab2),
  .a4b0(din_4_ab0), .a4b1(din_4_ab1),
  .a5b0(din_5_ab0), .a5b1(din_5_ab1),
  .a6b0(din_6_ab0),
  .a7b0(din_7_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_1_calc (
  .clk(clk), .p(addr_7_1),
  .a0b0(din_1_ab0), .a0b1(din_1_ab1), .a0b2(din_1_ab2), .a0b3(din_1_ab3),
  .a1b0(din_2_ab0), .a1b1(din_2_ab1), .a1b2(din_2_ab2), .a1b3(din_2_ab3),
  .a2b0(din_3_ab0), .a2b1(din_3_ab1), .a2b2(din_3_ab2),
  .a3b0(din_4_ab0), .a3b1(din_4_ab1), .a3b2(din_4_ab2),
  .a4b0(din_5_ab0), .a4b1(din_5_ab1),
  .a5b0(din_6_ab0), .a5b1(din_6_ab1),
  .a6b0(din_7_ab0),
  .a7b0(din_8_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_2_calc (
  .clk(clk), .p(addr_7_2),
  .a0b0(din_2_ab0), .a0b1(din_2_ab1), .a0b2(din_2_ab2), .a0b3(din_2_ab3),
  .a1b0(din_3_ab0), .a1b1(din_3_ab1), .a1b2(din_3_ab2), .a1b3(din_3_ab3),
  .a2b0(din_4_ab0), .a2b1(din_4_ab1), .a2b2(din_4_ab2),
  .a3b0(din_5_ab0), .a3b1(din_5_ab1), .a3b2(din_5_ab2),
  .a4b0(din_6_ab0), .a4b1(din_6_ab1),
  .a5b0(din_7_ab0), .a5b1(din_7_ab1),
  .a6b0(din_8_ab0),
  .a7b0(din_9_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_3_calc (
  .clk(clk), .p(addr_7_3),
  .a0b0(din_3_ab0), .a0b1(din_3_ab1), .a0b2(din_3_ab2), .a0b3(din_3_ab3),
  .a1b0(din_4_ab0), .a1b1(din_4_ab1), .a1b2(din_4_ab2), .a1b3(din_4_ab3),
  .a2b0(din_5_ab0), .a2b1(din_5_ab1), .a2b2(din_5_ab2),
  .a3b0(din_6_ab0), .a3b1(din_6_ab1), .a3b2(din_6_ab2),
  .a4b0(din_7_ab0), .a4b1(din_7_ab1),
  .a5b0(din_8_ab0), .a5b1(din_8_ab1),
  .a6b0(din_9_ab0),
  .a7b0(din_10_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_4_calc (
  .clk(clk), .p(addr_7_4),
  .a0b0(din_4_ab0), .a0b1(din_4_ab1), .a0b2(din_4_ab2), .a0b3(din_4_ab3),
  .a1b0(din_5_ab0), .a1b1(din_5_ab1), .a1b2(din_5_ab2), .a1b3(din_5_ab3),
  .a2b0(din_6_ab0), .a2b1(din_6_ab1), .a2b2(din_6_ab2),
  .a3b0(din_7_ab0), .a3b1(din_7_ab1), .a3b2(din_7_ab2),
  .a4b0(din_8_ab0), .a4b1(din_8_ab1),
  .a5b0(din_9_ab0), .a5b1(din_9_ab1),
  .a6b0(din_10_ab0),
  .a7b0(din_11_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_5_calc (
  .clk(clk), .p(addr_7_5),
  .a0b0(din_5_ab0), .a0b1(din_5_ab1), .a0b2(din_5_ab2), .a0b3(din_5_ab3),
  .a1b0(din_6_ab0), .a1b1(din_6_ab1), .a1b2(din_6_ab2), .a1b3(din_6_ab3),
  .a2b0(din_7_ab0), .a2b1(din_7_ab1), .a2b2(din_7_ab2),
  .a3b0(din_8_ab0), .a3b1(din_8_ab1), .a3b2(din_8_ab2),
  .a4b0(din_9_ab0), .a4b1(din_9_ab1),
  .a5b0(din_10_ab0), .a5b1(din_10_ab1),
  .a6b0(din_11_ab0),
  .a7b0(din_12_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_6_calc (
  .clk(clk), .p(addr_7_6),
  .a0b0(din_6_ab0), .a0b1(din_6_ab1), .a0b2(din_6_ab2), .a0b3(din_6_ab3),
  .a1b0(din_7_ab0), .a1b1(din_7_ab1), .a1b2(din_7_ab2), .a1b3(din_7_ab3),
  .a2b0(din_8_ab0), .a2b1(din_8_ab1), .a2b2(din_8_ab2),
  .a3b0(din_9_ab0), .a3b1(din_9_ab1), .a3b2(din_9_ab2),
  .a4b0(din_10_ab0), .a4b1(din_10_ab1),
  .a5b0(din_11_ab0), .a5b1(din_11_ab1),
  .a6b0(din_12_ab0),
  .a7b0(din_13_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_7_calc (
  .clk(clk), .p(addr_7_7),
  .a0b0(din_7_ab0), .a0b1(din_7_ab1), .a0b2(din_7_ab2), .a0b3(din_7_ab3),
  .a1b0(din_8_ab0), .a1b1(din_8_ab1), .a1b2(din_8_ab2), .a1b3(din_8_ab3),
  .a2b0(din_9_ab0), .a2b1(din_9_ab1), .a2b2(din_9_ab2),
  .a3b0(din_10_ab0), .a3b1(din_10_ab1), .a3b2(din_10_ab2),
  .a4b0(din_11_ab0), .a4b1(din_11_ab1),
  .a5b0(din_12_ab0), .a5b1(din_12_ab1),
  .a6b0(din_13_ab0),
  .a7b0(din_14_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_8_calc (
  .clk(clk), .p(addr_7_8),
  .a0b0(din_8_ab0), .a0b1(din_8_ab1), .a0b2(din_8_ab2), .a0b3(din_8_ab3),
  .a1b0(din_9_ab0), .a1b1(din_9_ab1), .a1b2(din_9_ab2), .a1b3(din_9_ab3),
  .a2b0(din_10_ab0), .a2b1(din_10_ab1), .a2b2(din_10_ab2),
  .a3b0(din_11_ab0), .a3b1(din_11_ab1), .a3b2(din_11_ab2),
  .a4b0(din_12_ab0), .a4b1(din_12_ab1),
  .a5b0(din_13_ab0), .a5b1(din_13_ab1),
  .a6b0(din_14_ab0),
  .a7b0(din_15_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_9_calc (
  .clk(clk), .p(addr_7_9),
  .a0b0(din_9_ab0), .a0b1(din_9_ab1), .a0b2(din_9_ab2), .a0b3(din_9_ab3),
  .a1b0(din_10_ab0), .a1b1(din_10_ab1), .a1b2(din_10_ab2), .a1b3(din_10_ab3),
  .a2b0(din_11_ab0), .a2b1(din_11_ab1), .a2b2(din_11_ab2),
  .a3b0(din_12_ab0), .a3b1(din_12_ab1), .a3b2(din_12_ab2),
  .a4b0(din_13_ab0), .a4b1(din_13_ab1),
  .a5b0(din_14_ab0), .a5b1(din_14_ab1),
  .a6b0(din_15_ab0),
  .a7b0(din_16_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_10_calc (
  .clk(clk), .p(addr_7_10),
  .a0b0(din_10_ab0), .a0b1(din_10_ab1), .a0b2(din_10_ab2), .a0b3(din_10_ab3),
  .a1b0(din_11_ab0), .a1b1(din_11_ab1), .a1b2(din_11_ab2), .a1b3(din_11_ab3),
  .a2b0(din_12_ab0), .a2b1(din_12_ab1), .a2b2(din_12_ab2),
  .a3b0(din_13_ab0), .a3b1(din_13_ab1), .a3b2(din_13_ab2),
  .a4b0(din_14_ab0), .a4b1(din_14_ab1),
  .a5b0(din_15_ab0), .a5b1(din_15_ab1),
  .a6b0(din_16_ab0),
  .a7b0(din_17_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_11_calc (
  .clk(clk), .p(addr_7_11),
  .a0b0(din_11_ab0), .a0b1(din_11_ab1), .a0b2(din_11_ab2), .a0b3(din_11_ab3),
  .a1b0(din_12_ab0), .a1b1(din_12_ab1), .a1b2(din_12_ab2), .a1b3(din_12_ab3),
  .a2b0(din_13_ab0), .a2b1(din_13_ab1), .a2b2(din_13_ab2),
  .a3b0(din_14_ab0), .a3b1(din_14_ab1), .a3b2(din_14_ab2),
  .a4b0(din_15_ab0), .a4b1(din_15_ab1),
  .a5b0(din_16_ab0), .a5b1(din_16_ab1),
  .a6b0(din_17_ab0),
  .a7b0(din_18_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_12_calc (
  .clk(clk), .p(addr_7_12),
  .a0b0(din_12_ab0), .a0b1(din_12_ab1), .a0b2(din_12_ab2), .a0b3(din_12_ab3),
  .a1b0(din_13_ab0), .a1b1(din_13_ab1), .a1b2(din_13_ab2), .a1b3(din_13_ab3),
  .a2b0(din_14_ab0), .a2b1(din_14_ab1), .a2b2(din_14_ab2),
  .a3b0(din_15_ab0), .a3b1(din_15_ab1), .a3b2(din_15_ab2),
  .a4b0(din_16_ab0), .a4b1(din_16_ab1),
  .a5b0(din_17_ab0), .a5b1(din_17_ab1),
  .a6b0(din_18_ab0),
  .a7b0(din_19_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_13_calc (
  .clk(clk), .p(addr_7_13),
  .a0b0(din_13_ab0), .a0b1(din_13_ab1), .a0b2(din_13_ab2), .a0b3(din_13_ab3),
  .a1b0(din_14_ab0), .a1b1(din_14_ab1), .a1b2(din_14_ab2), .a1b3(din_14_ab3),
  .a2b0(din_15_ab0), .a2b1(din_15_ab1), .a2b2(din_15_ab2),
  .a3b0(din_16_ab0), .a3b1(din_16_ab1), .a3b2(din_16_ab2),
  .a4b0(din_17_ab0), .a4b1(din_17_ab1),
  .a5b0(din_18_ab0), .a5b1(din_18_ab1),
  .a6b0(din_19_ab0),
  .a7b0(din_20_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_14_calc (
  .clk(clk), .p(addr_7_14),
  .a0b0(din_14_ab0), .a0b1(din_14_ab1), .a0b2(din_14_ab2), .a0b3(din_14_ab3),
  .a1b0(din_15_ab0), .a1b1(din_15_ab1), .a1b2(din_15_ab2), .a1b3(din_15_ab3),
  .a2b0(din_16_ab0), .a2b1(din_16_ab1), .a2b2(din_16_ab2),
  .a3b0(din_17_ab0), .a3b1(din_17_ab1), .a3b2(din_17_ab2),
  .a4b0(din_18_ab0), .a4b1(din_18_ab1),
  .a5b0(din_19_ab0), .a5b1(din_19_ab1),
  .a6b0(din_20_ab0),
  .a7b0(din_21_ab0)
);

acc_hash # (
	.ANDMSK(64'hff00000000000000),
	.NBITS(10)
) addr_7_15_calc (
  .clk(clk), .p(addr_7_15),
  .a0b0(din_15_ab0), .a0b1(din_15_ab1), .a0b2(din_15_ab2), .a0b3(din_15_ab3),
  .a1b0(din_16_ab0), .a1b1(din_16_ab1), .a1b2(din_16_ab2), .a1b3(din_16_ab3),
  .a2b0(din_17_ab0), .a2b1(din_17_ab1), .a2b2(din_17_ab2),
  .a3b0(din_18_ab0), .a3b1(din_18_ab1), .a3b2(din_18_ab2),
  .a4b0(din_19_ab0), .a4b1(din_19_ab1),
  .a5b0(din_20_ab0), .a5b1(din_20_ab1),
  .a6b0(din_21_ab0),
  .a7b0(din_22_ab0)
);




hashtable #(
    .NBITS(17),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(16384),
    .INIT_FILE("./src/memory_init/nf_bitmap0.mif")
)
hashtable_0_0 (
    .clk (clk),
	.addr0 (addr_0_0),
	.addr0_valid (addr_valid_0_0),
	.addr1 (addr_0_1),
	.addr1_valid (addr_valid_0_1),
    .dout0 (dout_0_0),
    .dout0_valid (dout_valid_0_0),
    .dout1 (dout_0_1),
    .dout1_valid (dout_valid_0_1)
);

hashtable #(
    .NBITS(17),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(16384),
    .INIT_FILE("./src/memory_init/nf_bitmap0.mif")
)
hashtable_0_1 (
    .clk (clk),
	.addr0 (addr_0_2),
	.addr0_valid (addr_valid_0_2),
	.addr1 (addr_0_3),
	.addr1_valid (addr_valid_0_3),
    .dout0 (dout_0_2),
    .dout0_valid (dout_valid_0_2),
    .dout1 (dout_0_3),
    .dout1_valid (dout_valid_0_3)
);

hashtable #(
    .NBITS(17),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(16384),
    .INIT_FILE("./src/memory_init/nf_bitmap0.mif")
)
hashtable_0_2 (
    .clk (clk),
	.addr0 (addr_0_4),
	.addr0_valid (addr_valid_0_4),
	.addr1 (addr_0_5),
	.addr1_valid (addr_valid_0_5),
    .dout0 (dout_0_4),
    .dout0_valid (dout_valid_0_4),
    .dout1 (dout_0_5),
    .dout1_valid (dout_valid_0_5)
);

hashtable #(
    .NBITS(17),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(16384),
    .INIT_FILE("./src/memory_init/nf_bitmap0.mif")
)
hashtable_0_3 (
    .clk (clk),
	.addr0 (addr_0_6),
	.addr0_valid (addr_valid_0_6),
	.addr1 (addr_0_7),
	.addr1_valid (addr_valid_0_7),
    .dout0 (dout_0_6),
    .dout0_valid (dout_valid_0_6),
    .dout1 (dout_0_7),
    .dout1_valid (dout_valid_0_7)
);

hashtable #(
    .NBITS(17),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(16384),
    .INIT_FILE("./src/memory_init/nf_bitmap0.mif")
)
hashtable_0_4 (
    .clk (clk),
	.addr0 (addr_0_8),
	.addr0_valid (addr_valid_0_8),
	.addr1 (addr_0_9),
	.addr1_valid (addr_valid_0_9),
    .dout0 (dout_0_8),
    .dout0_valid (dout_valid_0_8),
    .dout1 (dout_0_9),
    .dout1_valid (dout_valid_0_9)
);

hashtable #(
    .NBITS(17),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(16384),
    .INIT_FILE("./src/memory_init/nf_bitmap0.mif")
)
hashtable_0_5 (
    .clk (clk),
	.addr0 (addr_0_10),
	.addr0_valid (addr_valid_0_10),
	.addr1 (addr_0_11),
	.addr1_valid (addr_valid_0_11),
    .dout0 (dout_0_10),
    .dout0_valid (dout_valid_0_10),
    .dout1 (dout_0_11),
    .dout1_valid (dout_valid_0_11)
);

hashtable #(
    .NBITS(17),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(16384),
    .INIT_FILE("./src/memory_init/nf_bitmap0.mif")
)
hashtable_0_6 (
    .clk (clk),
	.addr0 (addr_0_12),
	.addr0_valid (addr_valid_0_12),
	.addr1 (addr_0_13),
	.addr1_valid (addr_valid_0_13),
    .dout0 (dout_0_12),
    .dout0_valid (dout_valid_0_12),
    .dout1 (dout_0_13),
    .dout1_valid (dout_valid_0_13)
);

hashtable #(
    .NBITS(17),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(16384),
    .INIT_FILE("./src/memory_init/nf_bitmap0.mif")
)
hashtable_0_7 (
    .clk (clk),
	.addr0 (addr_0_14),
	.addr0_valid (addr_valid_0_14),
	.addr1 (addr_0_15),
	.addr1_valid (addr_valid_0_15),
    .dout0 (dout_0_14),
    .dout0_valid (dout_valid_0_14),
    .dout1 (dout_0_15),
    .dout1_valid (dout_valid_0_15)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap1.mif")
)
hashtable_1_0 (
    .clk (clk),
	.addr0 (addr_1_0),
	.addr0_valid (addr_valid_1_0),
	.addr1 (addr_1_1),
	.addr1_valid (addr_valid_1_1),
    .dout0 (dout_1_0),
    .dout0_valid (dout_valid_1_0),
    .dout1 (dout_1_1),
    .dout1_valid (dout_valid_1_1)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap1.mif")
)
hashtable_1_1 (
    .clk (clk),
	.addr0 (addr_1_2),
	.addr0_valid (addr_valid_1_2),
	.addr1 (addr_1_3),
	.addr1_valid (addr_valid_1_3),
    .dout0 (dout_1_2),
    .dout0_valid (dout_valid_1_2),
    .dout1 (dout_1_3),
    .dout1_valid (dout_valid_1_3)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap1.mif")
)
hashtable_1_2 (
    .clk (clk),
	.addr0 (addr_1_4),
	.addr0_valid (addr_valid_1_4),
	.addr1 (addr_1_5),
	.addr1_valid (addr_valid_1_5),
    .dout0 (dout_1_4),
    .dout0_valid (dout_valid_1_4),
    .dout1 (dout_1_5),
    .dout1_valid (dout_valid_1_5)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap1.mif")
)
hashtable_1_3 (
    .clk (clk),
	.addr0 (addr_1_6),
	.addr0_valid (addr_valid_1_6),
	.addr1 (addr_1_7),
	.addr1_valid (addr_valid_1_7),
    .dout0 (dout_1_6),
    .dout0_valid (dout_valid_1_6),
    .dout1 (dout_1_7),
    .dout1_valid (dout_valid_1_7)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap1.mif")
)
hashtable_1_4 (
    .clk (clk),
	.addr0 (addr_1_8),
	.addr0_valid (addr_valid_1_8),
	.addr1 (addr_1_9),
	.addr1_valid (addr_valid_1_9),
    .dout0 (dout_1_8),
    .dout0_valid (dout_valid_1_8),
    .dout1 (dout_1_9),
    .dout1_valid (dout_valid_1_9)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap1.mif")
)
hashtable_1_5 (
    .clk (clk),
	.addr0 (addr_1_10),
	.addr0_valid (addr_valid_1_10),
	.addr1 (addr_1_11),
	.addr1_valid (addr_valid_1_11),
    .dout0 (dout_1_10),
    .dout0_valid (dout_valid_1_10),
    .dout1 (dout_1_11),
    .dout1_valid (dout_valid_1_11)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap1.mif")
)
hashtable_1_6 (
    .clk (clk),
	.addr0 (addr_1_12),
	.addr0_valid (addr_valid_1_12),
	.addr1 (addr_1_13),
	.addr1_valid (addr_valid_1_13),
    .dout0 (dout_1_12),
    .dout0_valid (dout_valid_1_12),
    .dout1 (dout_1_13),
    .dout1_valid (dout_valid_1_13)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap1.mif")
)
hashtable_1_7 (
    .clk (clk),
	.addr0 (addr_1_14),
	.addr0_valid (addr_valid_1_14),
	.addr1 (addr_1_15),
	.addr1_valid (addr_valid_1_15),
    .dout0 (dout_1_14),
    .dout0_valid (dout_valid_1_14),
    .dout1 (dout_1_15),
    .dout1_valid (dout_valid_1_15)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap2.mif")
)
hashtable_2_0 (
    .clk (clk),
	.addr0 (addr_2_0),
	.addr0_valid (addr_valid_2_0),
	.addr1 (addr_2_1),
	.addr1_valid (addr_valid_2_1),
    .dout0 (dout_2_0),
    .dout0_valid (dout_valid_2_0),
    .dout1 (dout_2_1),
    .dout1_valid (dout_valid_2_1)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap2.mif")
)
hashtable_2_1 (
    .clk (clk),
	.addr0 (addr_2_2),
	.addr0_valid (addr_valid_2_2),
	.addr1 (addr_2_3),
	.addr1_valid (addr_valid_2_3),
    .dout0 (dout_2_2),
    .dout0_valid (dout_valid_2_2),
    .dout1 (dout_2_3),
    .dout1_valid (dout_valid_2_3)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap2.mif")
)
hashtable_2_2 (
    .clk (clk),
	.addr0 (addr_2_4),
	.addr0_valid (addr_valid_2_4),
	.addr1 (addr_2_5),
	.addr1_valid (addr_valid_2_5),
    .dout0 (dout_2_4),
    .dout0_valid (dout_valid_2_4),
    .dout1 (dout_2_5),
    .dout1_valid (dout_valid_2_5)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap2.mif")
)
hashtable_2_3 (
    .clk (clk),
	.addr0 (addr_2_6),
	.addr0_valid (addr_valid_2_6),
	.addr1 (addr_2_7),
	.addr1_valid (addr_valid_2_7),
    .dout0 (dout_2_6),
    .dout0_valid (dout_valid_2_6),
    .dout1 (dout_2_7),
    .dout1_valid (dout_valid_2_7)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap2.mif")
)
hashtable_2_4 (
    .clk (clk),
	.addr0 (addr_2_8),
	.addr0_valid (addr_valid_2_8),
	.addr1 (addr_2_9),
	.addr1_valid (addr_valid_2_9),
    .dout0 (dout_2_8),
    .dout0_valid (dout_valid_2_8),
    .dout1 (dout_2_9),
    .dout1_valid (dout_valid_2_9)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap2.mif")
)
hashtable_2_5 (
    .clk (clk),
	.addr0 (addr_2_10),
	.addr0_valid (addr_valid_2_10),
	.addr1 (addr_2_11),
	.addr1_valid (addr_valid_2_11),
    .dout0 (dout_2_10),
    .dout0_valid (dout_valid_2_10),
    .dout1 (dout_2_11),
    .dout1_valid (dout_valid_2_11)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap2.mif")
)
hashtable_2_6 (
    .clk (clk),
	.addr0 (addr_2_12),
	.addr0_valid (addr_valid_2_12),
	.addr1 (addr_2_13),
	.addr1_valid (addr_valid_2_13),
    .dout0 (dout_2_12),
    .dout0_valid (dout_valid_2_12),
    .dout1 (dout_2_13),
    .dout1_valid (dout_valid_2_13)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap2.mif")
)
hashtable_2_7 (
    .clk (clk),
	.addr0 (addr_2_14),
	.addr0_valid (addr_valid_2_14),
	.addr1 (addr_2_15),
	.addr1_valid (addr_valid_2_15),
    .dout0 (dout_2_14),
    .dout0_valid (dout_valid_2_14),
    .dout1 (dout_2_15),
    .dout1_valid (dout_valid_2_15)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap3.mif")
)
hashtable_3_0 (
    .clk (clk),
	.addr0 (addr_3_0),
	.addr0_valid (addr_valid_3_0),
	.addr1 (addr_3_1),
	.addr1_valid (addr_valid_3_1),
    .dout0 (dout_3_0),
    .dout0_valid (dout_valid_3_0),
    .dout1 (dout_3_1),
    .dout1_valid (dout_valid_3_1)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap3.mif")
)
hashtable_3_1 (
    .clk (clk),
	.addr0 (addr_3_2),
	.addr0_valid (addr_valid_3_2),
	.addr1 (addr_3_3),
	.addr1_valid (addr_valid_3_3),
    .dout0 (dout_3_2),
    .dout0_valid (dout_valid_3_2),
    .dout1 (dout_3_3),
    .dout1_valid (dout_valid_3_3)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap3.mif")
)
hashtable_3_2 (
    .clk (clk),
	.addr0 (addr_3_4),
	.addr0_valid (addr_valid_3_4),
	.addr1 (addr_3_5),
	.addr1_valid (addr_valid_3_5),
    .dout0 (dout_3_4),
    .dout0_valid (dout_valid_3_4),
    .dout1 (dout_3_5),
    .dout1_valid (dout_valid_3_5)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap3.mif")
)
hashtable_3_3 (
    .clk (clk),
	.addr0 (addr_3_6),
	.addr0_valid (addr_valid_3_6),
	.addr1 (addr_3_7),
	.addr1_valid (addr_valid_3_7),
    .dout0 (dout_3_6),
    .dout0_valid (dout_valid_3_6),
    .dout1 (dout_3_7),
    .dout1_valid (dout_valid_3_7)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap3.mif")
)
hashtable_3_4 (
    .clk (clk),
	.addr0 (addr_3_8),
	.addr0_valid (addr_valid_3_8),
	.addr1 (addr_3_9),
	.addr1_valid (addr_valid_3_9),
    .dout0 (dout_3_8),
    .dout0_valid (dout_valid_3_8),
    .dout1 (dout_3_9),
    .dout1_valid (dout_valid_3_9)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap3.mif")
)
hashtable_3_5 (
    .clk (clk),
	.addr0 (addr_3_10),
	.addr0_valid (addr_valid_3_10),
	.addr1 (addr_3_11),
	.addr1_valid (addr_valid_3_11),
    .dout0 (dout_3_10),
    .dout0_valid (dout_valid_3_10),
    .dout1 (dout_3_11),
    .dout1_valid (dout_valid_3_11)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap3.mif")
)
hashtable_3_6 (
    .clk (clk),
	.addr0 (addr_3_12),
	.addr0_valid (addr_valid_3_12),
	.addr1 (addr_3_13),
	.addr1_valid (addr_valid_3_13),
    .dout0 (dout_3_12),
    .dout0_valid (dout_valid_3_12),
    .dout1 (dout_3_13),
    .dout1_valid (dout_valid_3_13)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap3.mif")
)
hashtable_3_7 (
    .clk (clk),
	.addr0 (addr_3_14),
	.addr0_valid (addr_valid_3_14),
	.addr1 (addr_3_15),
	.addr1_valid (addr_valid_3_15),
    .dout0 (dout_3_14),
    .dout0_valid (dout_valid_3_14),
    .dout1 (dout_3_15),
    .dout1_valid (dout_valid_3_15)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap4.mif")
)
hashtable_4_0 (
    .clk (clk),
	.addr0 (addr_4_0),
	.addr0_valid (addr_valid_4_0),
	.addr1 (addr_4_1),
	.addr1_valid (addr_valid_4_1),
    .dout0 (dout_4_0),
    .dout0_valid (dout_valid_4_0),
    .dout1 (dout_4_1),
    .dout1_valid (dout_valid_4_1)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap4.mif")
)
hashtable_4_1 (
    .clk (clk),
	.addr0 (addr_4_2),
	.addr0_valid (addr_valid_4_2),
	.addr1 (addr_4_3),
	.addr1_valid (addr_valid_4_3),
    .dout0 (dout_4_2),
    .dout0_valid (dout_valid_4_2),
    .dout1 (dout_4_3),
    .dout1_valid (dout_valid_4_3)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap4.mif")
)
hashtable_4_2 (
    .clk (clk),
	.addr0 (addr_4_4),
	.addr0_valid (addr_valid_4_4),
	.addr1 (addr_4_5),
	.addr1_valid (addr_valid_4_5),
    .dout0 (dout_4_4),
    .dout0_valid (dout_valid_4_4),
    .dout1 (dout_4_5),
    .dout1_valid (dout_valid_4_5)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap4.mif")
)
hashtable_4_3 (
    .clk (clk),
	.addr0 (addr_4_6),
	.addr0_valid (addr_valid_4_6),
	.addr1 (addr_4_7),
	.addr1_valid (addr_valid_4_7),
    .dout0 (dout_4_6),
    .dout0_valid (dout_valid_4_6),
    .dout1 (dout_4_7),
    .dout1_valid (dout_valid_4_7)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap4.mif")
)
hashtable_4_4 (
    .clk (clk),
	.addr0 (addr_4_8),
	.addr0_valid (addr_valid_4_8),
	.addr1 (addr_4_9),
	.addr1_valid (addr_valid_4_9),
    .dout0 (dout_4_8),
    .dout0_valid (dout_valid_4_8),
    .dout1 (dout_4_9),
    .dout1_valid (dout_valid_4_9)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap4.mif")
)
hashtable_4_5 (
    .clk (clk),
	.addr0 (addr_4_10),
	.addr0_valid (addr_valid_4_10),
	.addr1 (addr_4_11),
	.addr1_valid (addr_valid_4_11),
    .dout0 (dout_4_10),
    .dout0_valid (dout_valid_4_10),
    .dout1 (dout_4_11),
    .dout1_valid (dout_valid_4_11)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap4.mif")
)
hashtable_4_6 (
    .clk (clk),
	.addr0 (addr_4_12),
	.addr0_valid (addr_valid_4_12),
	.addr1 (addr_4_13),
	.addr1_valid (addr_valid_4_13),
    .dout0 (dout_4_12),
    .dout0_valid (dout_valid_4_12),
    .dout1 (dout_4_13),
    .dout1_valid (dout_valid_4_13)
);

hashtable #(
    .NBITS(13),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(1024),
    .INIT_FILE("./src/memory_init/nf_bitmap4.mif")
)
hashtable_4_7 (
    .clk (clk),
	.addr0 (addr_4_14),
	.addr0_valid (addr_valid_4_14),
	.addr1 (addr_4_15),
	.addr1_valid (addr_valid_4_15),
    .dout0 (dout_4_14),
    .dout0_valid (dout_valid_4_14),
    .dout1 (dout_4_15),
    .dout1_valid (dout_valid_4_15)
);

hashtable #(
    .NBITS(12),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(512),
    .INIT_FILE("./src/memory_init/nf_bitmap5.mif")
)
hashtable_5_0 (
    .clk (clk),
	.addr0 (addr_5_0),
	.addr0_valid (addr_valid_5_0),
	.addr1 (addr_5_1),
	.addr1_valid (addr_valid_5_1),
    .dout0 (dout_5_0),
    .dout0_valid (dout_valid_5_0),
    .dout1 (dout_5_1),
    .dout1_valid (dout_valid_5_1)
);

hashtable #(
    .NBITS(12),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(512),
    .INIT_FILE("./src/memory_init/nf_bitmap5.mif")
)
hashtable_5_1 (
    .clk (clk),
	.addr0 (addr_5_2),
	.addr0_valid (addr_valid_5_2),
	.addr1 (addr_5_3),
	.addr1_valid (addr_valid_5_3),
    .dout0 (dout_5_2),
    .dout0_valid (dout_valid_5_2),
    .dout1 (dout_5_3),
    .dout1_valid (dout_valid_5_3)
);

hashtable #(
    .NBITS(12),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(512),
    .INIT_FILE("./src/memory_init/nf_bitmap5.mif")
)
hashtable_5_2 (
    .clk (clk),
	.addr0 (addr_5_4),
	.addr0_valid (addr_valid_5_4),
	.addr1 (addr_5_5),
	.addr1_valid (addr_valid_5_5),
    .dout0 (dout_5_4),
    .dout0_valid (dout_valid_5_4),
    .dout1 (dout_5_5),
    .dout1_valid (dout_valid_5_5)
);

hashtable #(
    .NBITS(12),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(512),
    .INIT_FILE("./src/memory_init/nf_bitmap5.mif")
)
hashtable_5_3 (
    .clk (clk),
	.addr0 (addr_5_6),
	.addr0_valid (addr_valid_5_6),
	.addr1 (addr_5_7),
	.addr1_valid (addr_valid_5_7),
    .dout0 (dout_5_6),
    .dout0_valid (dout_valid_5_6),
    .dout1 (dout_5_7),
    .dout1_valid (dout_valid_5_7)
);

hashtable #(
    .NBITS(12),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(512),
    .INIT_FILE("./src/memory_init/nf_bitmap5.mif")
)
hashtable_5_4 (
    .clk (clk),
	.addr0 (addr_5_8),
	.addr0_valid (addr_valid_5_8),
	.addr1 (addr_5_9),
	.addr1_valid (addr_valid_5_9),
    .dout0 (dout_5_8),
    .dout0_valid (dout_valid_5_8),
    .dout1 (dout_5_9),
    .dout1_valid (dout_valid_5_9)
);

hashtable #(
    .NBITS(12),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(512),
    .INIT_FILE("./src/memory_init/nf_bitmap5.mif")
)
hashtable_5_5 (
    .clk (clk),
	.addr0 (addr_5_10),
	.addr0_valid (addr_valid_5_10),
	.addr1 (addr_5_11),
	.addr1_valid (addr_valid_5_11),
    .dout0 (dout_5_10),
    .dout0_valid (dout_valid_5_10),
    .dout1 (dout_5_11),
    .dout1_valid (dout_valid_5_11)
);

hashtable #(
    .NBITS(12),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(512),
    .INIT_FILE("./src/memory_init/nf_bitmap5.mif")
)
hashtable_5_6 (
    .clk (clk),
	.addr0 (addr_5_12),
	.addr0_valid (addr_valid_5_12),
	.addr1 (addr_5_13),
	.addr1_valid (addr_valid_5_13),
    .dout0 (dout_5_12),
    .dout0_valid (dout_valid_5_12),
    .dout1 (dout_5_13),
    .dout1_valid (dout_valid_5_13)
);

hashtable #(
    .NBITS(12),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(512),
    .INIT_FILE("./src/memory_init/nf_bitmap5.mif")
)
hashtable_5_7 (
    .clk (clk),
	.addr0 (addr_5_14),
	.addr0_valid (addr_valid_5_14),
	.addr1 (addr_5_15),
	.addr1_valid (addr_valid_5_15),
    .dout0 (dout_5_14),
    .dout0_valid (dout_valid_5_14),
    .dout1 (dout_5_15),
    .dout1_valid (dout_valid_5_15)
);

hashtable #(
    .NBITS(11),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(256),
    .INIT_FILE("./src/memory_init/nf_bitmap6.mif")
)
hashtable_6_0 (
    .clk (clk),
	.addr0 (addr_6_0),
	.addr0_valid (addr_valid_6_0),
	.addr1 (addr_6_1),
	.addr1_valid (addr_valid_6_1),
    .dout0 (dout_6_0),
    .dout0_valid (dout_valid_6_0),
    .dout1 (dout_6_1),
    .dout1_valid (dout_valid_6_1)
);

hashtable #(
    .NBITS(11),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(256),
    .INIT_FILE("./src/memory_init/nf_bitmap6.mif")
)
hashtable_6_1 (
    .clk (clk),
	.addr0 (addr_6_2),
	.addr0_valid (addr_valid_6_2),
	.addr1 (addr_6_3),
	.addr1_valid (addr_valid_6_3),
    .dout0 (dout_6_2),
    .dout0_valid (dout_valid_6_2),
    .dout1 (dout_6_3),
    .dout1_valid (dout_valid_6_3)
);

hashtable #(
    .NBITS(11),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(256),
    .INIT_FILE("./src/memory_init/nf_bitmap6.mif")
)
hashtable_6_2 (
    .clk (clk),
	.addr0 (addr_6_4),
	.addr0_valid (addr_valid_6_4),
	.addr1 (addr_6_5),
	.addr1_valid (addr_valid_6_5),
    .dout0 (dout_6_4),
    .dout0_valid (dout_valid_6_4),
    .dout1 (dout_6_5),
    .dout1_valid (dout_valid_6_5)
);

hashtable #(
    .NBITS(11),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(256),
    .INIT_FILE("./src/memory_init/nf_bitmap6.mif")
)
hashtable_6_3 (
    .clk (clk),
	.addr0 (addr_6_6),
	.addr0_valid (addr_valid_6_6),
	.addr1 (addr_6_7),
	.addr1_valid (addr_valid_6_7),
    .dout0 (dout_6_6),
    .dout0_valid (dout_valid_6_6),
    .dout1 (dout_6_7),
    .dout1_valid (dout_valid_6_7)
);

hashtable #(
    .NBITS(11),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(256),
    .INIT_FILE("./src/memory_init/nf_bitmap6.mif")
)
hashtable_6_4 (
    .clk (clk),
	.addr0 (addr_6_8),
	.addr0_valid (addr_valid_6_8),
	.addr1 (addr_6_9),
	.addr1_valid (addr_valid_6_9),
    .dout0 (dout_6_8),
    .dout0_valid (dout_valid_6_8),
    .dout1 (dout_6_9),
    .dout1_valid (dout_valid_6_9)
);

hashtable #(
    .NBITS(11),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(256),
    .INIT_FILE("./src/memory_init/nf_bitmap6.mif")
)
hashtable_6_5 (
    .clk (clk),
	.addr0 (addr_6_10),
	.addr0_valid (addr_valid_6_10),
	.addr1 (addr_6_11),
	.addr1_valid (addr_valid_6_11),
    .dout0 (dout_6_10),
    .dout0_valid (dout_valid_6_10),
    .dout1 (dout_6_11),
    .dout1_valid (dout_valid_6_11)
);

hashtable #(
    .NBITS(11),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(256),
    .INIT_FILE("./src/memory_init/nf_bitmap6.mif")
)
hashtable_6_6 (
    .clk (clk),
	.addr0 (addr_6_12),
	.addr0_valid (addr_valid_6_12),
	.addr1 (addr_6_13),
	.addr1_valid (addr_valid_6_13),
    .dout0 (dout_6_12),
    .dout0_valid (dout_valid_6_12),
    .dout1 (dout_6_13),
    .dout1_valid (dout_valid_6_13)
);

hashtable #(
    .NBITS(11),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(256),
    .INIT_FILE("./src/memory_init/nf_bitmap6.mif")
)
hashtable_6_7 (
    .clk (clk),
	.addr0 (addr_6_14),
	.addr0_valid (addr_valid_6_14),
	.addr1 (addr_6_15),
	.addr1_valid (addr_valid_6_15),
    .dout0 (dout_6_14),
    .dout0_valid (dout_valid_6_14),
    .dout1 (dout_6_15),
    .dout1_valid (dout_valid_6_15)
);

hashtable #(
    .NBITS(10),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(128),
    .INIT_FILE("./src/memory_init/nf_bitmap7.mif")
)
hashtable_7_0 (
    .clk (clk),
	.addr0 (addr_7_0),
	.addr0_valid (addr_valid_7_0),
	.addr1 (addr_7_1),
	.addr1_valid (addr_valid_7_1),
    .dout0 (dout_7_0),
    .dout0_valid (dout_valid_7_0),
    .dout1 (dout_7_1),
    .dout1_valid (dout_valid_7_1)
);

hashtable #(
    .NBITS(10),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(128),
    .INIT_FILE("./src/memory_init/nf_bitmap7.mif")
)
hashtable_7_1 (
    .clk (clk),
	.addr0 (addr_7_2),
	.addr0_valid (addr_valid_7_2),
	.addr1 (addr_7_3),
	.addr1_valid (addr_valid_7_3),
    .dout0 (dout_7_2),
    .dout0_valid (dout_valid_7_2),
    .dout1 (dout_7_3),
    .dout1_valid (dout_valid_7_3)
);

hashtable #(
    .NBITS(10),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(128),
    .INIT_FILE("./src/memory_init/nf_bitmap7.mif")
)
hashtable_7_2 (
    .clk (clk),
	.addr0 (addr_7_4),
	.addr0_valid (addr_valid_7_4),
	.addr1 (addr_7_5),
	.addr1_valid (addr_valid_7_5),
    .dout0 (dout_7_4),
    .dout0_valid (dout_valid_7_4),
    .dout1 (dout_7_5),
    .dout1_valid (dout_valid_7_5)
);

hashtable #(
    .NBITS(10),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(128),
    .INIT_FILE("./src/memory_init/nf_bitmap7.mif")
)
hashtable_7_3 (
    .clk (clk),
	.addr0 (addr_7_6),
	.addr0_valid (addr_valid_7_6),
	.addr1 (addr_7_7),
	.addr1_valid (addr_valid_7_7),
    .dout0 (dout_7_6),
    .dout0_valid (dout_valid_7_6),
    .dout1 (dout_7_7),
    .dout1_valid (dout_valid_7_7)
);

hashtable #(
    .NBITS(10),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(128),
    .INIT_FILE("./src/memory_init/nf_bitmap7.mif")
)
hashtable_7_4 (
    .clk (clk),
	.addr0 (addr_7_8),
	.addr0_valid (addr_valid_7_8),
	.addr1 (addr_7_9),
	.addr1_valid (addr_valid_7_9),
    .dout0 (dout_7_8),
    .dout0_valid (dout_valid_7_8),
    .dout1 (dout_7_9),
    .dout1_valid (dout_valid_7_9)
);

hashtable #(
    .NBITS(10),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(128),
    .INIT_FILE("./src/memory_init/nf_bitmap7.mif")
)
hashtable_7_5 (
    .clk (clk),
	.addr0 (addr_7_10),
	.addr0_valid (addr_valid_7_10),
	.addr1 (addr_7_11),
	.addr1_valid (addr_valid_7_11),
    .dout0 (dout_7_10),
    .dout0_valid (dout_valid_7_10),
    .dout1 (dout_7_11),
    .dout1_valid (dout_valid_7_11)
);

hashtable #(
    .NBITS(10),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(128),
    .INIT_FILE("./src/memory_init/nf_bitmap7.mif")
)
hashtable_7_6 (
    .clk (clk),
	.addr0 (addr_7_12),
	.addr0_valid (addr_valid_7_12),
	.addr1 (addr_7_13),
	.addr1_valid (addr_valid_7_13),
    .dout0 (dout_7_12),
    .dout0_valid (dout_valid_7_12),
    .dout1 (dout_7_13),
    .dout1_valid (dout_valid_7_13)
);

hashtable #(
    .NBITS(10),
    .DWIDTH(NF_WIDTH),
    .MEM_SIZE(128),
    .INIT_FILE("./src/memory_init/nf_bitmap7.mif")
)
hashtable_7_7 (
    .clk (clk),
	.addr0 (addr_7_14),
	.addr0_valid (addr_valid_7_14),
	.addr1 (addr_7_15),
	.addr1_valid (addr_valid_7_15),
    .dout0 (dout_7_14),
    .dout0_valid (dout_valid_7_14),
    .dout1 (dout_7_15),
    .dout1_valid (dout_valid_7_15)
);

endmodule
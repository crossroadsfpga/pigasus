`include "./src/struct_s.sv"
//`define DUMMY
module frontend (clk,rst,
    hash_out_0_0,
    hash_out_valid_filter_0_0,
    hash_out_0_1,
    hash_out_valid_filter_0_1,
    hash_out_0_2,
    hash_out_valid_filter_0_2,
    hash_out_0_3,
    hash_out_valid_filter_0_3,
    hash_out_0_4,
    hash_out_valid_filter_0_4,
    hash_out_0_5,
    hash_out_valid_filter_0_5,
    hash_out_0_6,
    hash_out_valid_filter_0_6,
    hash_out_0_7,
    hash_out_valid_filter_0_7,
    hash_out_0_8,
    hash_out_valid_filter_0_8,
    hash_out_0_9,
    hash_out_valid_filter_0_9,
    hash_out_0_10,
    hash_out_valid_filter_0_10,
    hash_out_0_11,
    hash_out_valid_filter_0_11,
    hash_out_0_12,
    hash_out_valid_filter_0_12,
    hash_out_0_13,
    hash_out_valid_filter_0_13,
    hash_out_0_14,
    hash_out_valid_filter_0_14,
    hash_out_0_15,
    hash_out_valid_filter_0_15,
    hash_out_0_16,
    hash_out_valid_filter_0_16,
    hash_out_0_17,
    hash_out_valid_filter_0_17,
    hash_out_0_18,
    hash_out_valid_filter_0_18,
    hash_out_0_19,
    hash_out_valid_filter_0_19,
    hash_out_0_20,
    hash_out_valid_filter_0_20,
    hash_out_0_21,
    hash_out_valid_filter_0_21,
    hash_out_0_22,
    hash_out_valid_filter_0_22,
    hash_out_0_23,
    hash_out_valid_filter_0_23,
    hash_out_0_24,
    hash_out_valid_filter_0_24,
    hash_out_0_25,
    hash_out_valid_filter_0_25,
    hash_out_0_26,
    hash_out_valid_filter_0_26,
    hash_out_0_27,
    hash_out_valid_filter_0_27,
    hash_out_0_28,
    hash_out_valid_filter_0_28,
    hash_out_0_29,
    hash_out_valid_filter_0_29,
    hash_out_0_30,
    hash_out_valid_filter_0_30,
    hash_out_0_31,
    hash_out_valid_filter_0_31,
    hash_out_1_0,
    hash_out_valid_filter_1_0,
    hash_out_1_1,
    hash_out_valid_filter_1_1,
    hash_out_1_2,
    hash_out_valid_filter_1_2,
    hash_out_1_3,
    hash_out_valid_filter_1_3,
    hash_out_1_4,
    hash_out_valid_filter_1_4,
    hash_out_1_5,
    hash_out_valid_filter_1_5,
    hash_out_1_6,
    hash_out_valid_filter_1_6,
    hash_out_1_7,
    hash_out_valid_filter_1_7,
    hash_out_1_8,
    hash_out_valid_filter_1_8,
    hash_out_1_9,
    hash_out_valid_filter_1_9,
    hash_out_1_10,
    hash_out_valid_filter_1_10,
    hash_out_1_11,
    hash_out_valid_filter_1_11,
    hash_out_1_12,
    hash_out_valid_filter_1_12,
    hash_out_1_13,
    hash_out_valid_filter_1_13,
    hash_out_1_14,
    hash_out_valid_filter_1_14,
    hash_out_1_15,
    hash_out_valid_filter_1_15,
    hash_out_1_16,
    hash_out_valid_filter_1_16,
    hash_out_1_17,
    hash_out_valid_filter_1_17,
    hash_out_1_18,
    hash_out_valid_filter_1_18,
    hash_out_1_19,
    hash_out_valid_filter_1_19,
    hash_out_1_20,
    hash_out_valid_filter_1_20,
    hash_out_1_21,
    hash_out_valid_filter_1_21,
    hash_out_1_22,
    hash_out_valid_filter_1_22,
    hash_out_1_23,
    hash_out_valid_filter_1_23,
    hash_out_1_24,
    hash_out_valid_filter_1_24,
    hash_out_1_25,
    hash_out_valid_filter_1_25,
    hash_out_1_26,
    hash_out_valid_filter_1_26,
    hash_out_1_27,
    hash_out_valid_filter_1_27,
    hash_out_1_28,
    hash_out_valid_filter_1_28,
    hash_out_1_29,
    hash_out_valid_filter_1_29,
    hash_out_1_30,
    hash_out_valid_filter_1_30,
    hash_out_1_31,
    hash_out_valid_filter_1_31,
    hash_out_2_0,
    hash_out_valid_filter_2_0,
    hash_out_2_1,
    hash_out_valid_filter_2_1,
    hash_out_2_2,
    hash_out_valid_filter_2_2,
    hash_out_2_3,
    hash_out_valid_filter_2_3,
    hash_out_2_4,
    hash_out_valid_filter_2_4,
    hash_out_2_5,
    hash_out_valid_filter_2_5,
    hash_out_2_6,
    hash_out_valid_filter_2_6,
    hash_out_2_7,
    hash_out_valid_filter_2_7,
    hash_out_2_8,
    hash_out_valid_filter_2_8,
    hash_out_2_9,
    hash_out_valid_filter_2_9,
    hash_out_2_10,
    hash_out_valid_filter_2_10,
    hash_out_2_11,
    hash_out_valid_filter_2_11,
    hash_out_2_12,
    hash_out_valid_filter_2_12,
    hash_out_2_13,
    hash_out_valid_filter_2_13,
    hash_out_2_14,
    hash_out_valid_filter_2_14,
    hash_out_2_15,
    hash_out_valid_filter_2_15,
    hash_out_2_16,
    hash_out_valid_filter_2_16,
    hash_out_2_17,
    hash_out_valid_filter_2_17,
    hash_out_2_18,
    hash_out_valid_filter_2_18,
    hash_out_2_19,
    hash_out_valid_filter_2_19,
    hash_out_2_20,
    hash_out_valid_filter_2_20,
    hash_out_2_21,
    hash_out_valid_filter_2_21,
    hash_out_2_22,
    hash_out_valid_filter_2_22,
    hash_out_2_23,
    hash_out_valid_filter_2_23,
    hash_out_2_24,
    hash_out_valid_filter_2_24,
    hash_out_2_25,
    hash_out_valid_filter_2_25,
    hash_out_2_26,
    hash_out_valid_filter_2_26,
    hash_out_2_27,
    hash_out_valid_filter_2_27,
    hash_out_2_28,
    hash_out_valid_filter_2_28,
    hash_out_2_29,
    hash_out_valid_filter_2_29,
    hash_out_2_30,
    hash_out_valid_filter_2_30,
    hash_out_2_31,
    hash_out_valid_filter_2_31,
    hash_out_3_0,
    hash_out_valid_filter_3_0,
    hash_out_3_1,
    hash_out_valid_filter_3_1,
    hash_out_3_2,
    hash_out_valid_filter_3_2,
    hash_out_3_3,
    hash_out_valid_filter_3_3,
    hash_out_3_4,
    hash_out_valid_filter_3_4,
    hash_out_3_5,
    hash_out_valid_filter_3_5,
    hash_out_3_6,
    hash_out_valid_filter_3_6,
    hash_out_3_7,
    hash_out_valid_filter_3_7,
    hash_out_3_8,
    hash_out_valid_filter_3_8,
    hash_out_3_9,
    hash_out_valid_filter_3_9,
    hash_out_3_10,
    hash_out_valid_filter_3_10,
    hash_out_3_11,
    hash_out_valid_filter_3_11,
    hash_out_3_12,
    hash_out_valid_filter_3_12,
    hash_out_3_13,
    hash_out_valid_filter_3_13,
    hash_out_3_14,
    hash_out_valid_filter_3_14,
    hash_out_3_15,
    hash_out_valid_filter_3_15,
    hash_out_3_16,
    hash_out_valid_filter_3_16,
    hash_out_3_17,
    hash_out_valid_filter_3_17,
    hash_out_3_18,
    hash_out_valid_filter_3_18,
    hash_out_3_19,
    hash_out_valid_filter_3_19,
    hash_out_3_20,
    hash_out_valid_filter_3_20,
    hash_out_3_21,
    hash_out_valid_filter_3_21,
    hash_out_3_22,
    hash_out_valid_filter_3_22,
    hash_out_3_23,
    hash_out_valid_filter_3_23,
    hash_out_3_24,
    hash_out_valid_filter_3_24,
    hash_out_3_25,
    hash_out_valid_filter_3_25,
    hash_out_3_26,
    hash_out_valid_filter_3_26,
    hash_out_3_27,
    hash_out_valid_filter_3_27,
    hash_out_3_28,
    hash_out_valid_filter_3_28,
    hash_out_3_29,
    hash_out_valid_filter_3_29,
    hash_out_3_30,
    hash_out_valid_filter_3_30,
    hash_out_3_31,
    hash_out_valid_filter_3_31,
    hash_out_4_0,
    hash_out_valid_filter_4_0,
    hash_out_4_1,
    hash_out_valid_filter_4_1,
    hash_out_4_2,
    hash_out_valid_filter_4_2,
    hash_out_4_3,
    hash_out_valid_filter_4_3,
    hash_out_4_4,
    hash_out_valid_filter_4_4,
    hash_out_4_5,
    hash_out_valid_filter_4_5,
    hash_out_4_6,
    hash_out_valid_filter_4_6,
    hash_out_4_7,
    hash_out_valid_filter_4_7,
    hash_out_4_8,
    hash_out_valid_filter_4_8,
    hash_out_4_9,
    hash_out_valid_filter_4_9,
    hash_out_4_10,
    hash_out_valid_filter_4_10,
    hash_out_4_11,
    hash_out_valid_filter_4_11,
    hash_out_4_12,
    hash_out_valid_filter_4_12,
    hash_out_4_13,
    hash_out_valid_filter_4_13,
    hash_out_4_14,
    hash_out_valid_filter_4_14,
    hash_out_4_15,
    hash_out_valid_filter_4_15,
    hash_out_4_16,
    hash_out_valid_filter_4_16,
    hash_out_4_17,
    hash_out_valid_filter_4_17,
    hash_out_4_18,
    hash_out_valid_filter_4_18,
    hash_out_4_19,
    hash_out_valid_filter_4_19,
    hash_out_4_20,
    hash_out_valid_filter_4_20,
    hash_out_4_21,
    hash_out_valid_filter_4_21,
    hash_out_4_22,
    hash_out_valid_filter_4_22,
    hash_out_4_23,
    hash_out_valid_filter_4_23,
    hash_out_4_24,
    hash_out_valid_filter_4_24,
    hash_out_4_25,
    hash_out_valid_filter_4_25,
    hash_out_4_26,
    hash_out_valid_filter_4_26,
    hash_out_4_27,
    hash_out_valid_filter_4_27,
    hash_out_4_28,
    hash_out_valid_filter_4_28,
    hash_out_4_29,
    hash_out_valid_filter_4_29,
    hash_out_4_30,
    hash_out_valid_filter_4_30,
    hash_out_4_31,
    hash_out_valid_filter_4_31,
    hash_out_5_0,
    hash_out_valid_filter_5_0,
    hash_out_5_1,
    hash_out_valid_filter_5_1,
    hash_out_5_2,
    hash_out_valid_filter_5_2,
    hash_out_5_3,
    hash_out_valid_filter_5_3,
    hash_out_5_4,
    hash_out_valid_filter_5_4,
    hash_out_5_5,
    hash_out_valid_filter_5_5,
    hash_out_5_6,
    hash_out_valid_filter_5_6,
    hash_out_5_7,
    hash_out_valid_filter_5_7,
    hash_out_5_8,
    hash_out_valid_filter_5_8,
    hash_out_5_9,
    hash_out_valid_filter_5_9,
    hash_out_5_10,
    hash_out_valid_filter_5_10,
    hash_out_5_11,
    hash_out_valid_filter_5_11,
    hash_out_5_12,
    hash_out_valid_filter_5_12,
    hash_out_5_13,
    hash_out_valid_filter_5_13,
    hash_out_5_14,
    hash_out_valid_filter_5_14,
    hash_out_5_15,
    hash_out_valid_filter_5_15,
    hash_out_5_16,
    hash_out_valid_filter_5_16,
    hash_out_5_17,
    hash_out_valid_filter_5_17,
    hash_out_5_18,
    hash_out_valid_filter_5_18,
    hash_out_5_19,
    hash_out_valid_filter_5_19,
    hash_out_5_20,
    hash_out_valid_filter_5_20,
    hash_out_5_21,
    hash_out_valid_filter_5_21,
    hash_out_5_22,
    hash_out_valid_filter_5_22,
    hash_out_5_23,
    hash_out_valid_filter_5_23,
    hash_out_5_24,
    hash_out_valid_filter_5_24,
    hash_out_5_25,
    hash_out_valid_filter_5_25,
    hash_out_5_26,
    hash_out_valid_filter_5_26,
    hash_out_5_27,
    hash_out_valid_filter_5_27,
    hash_out_5_28,
    hash_out_valid_filter_5_28,
    hash_out_5_29,
    hash_out_valid_filter_5_29,
    hash_out_5_30,
    hash_out_valid_filter_5_30,
    hash_out_5_31,
    hash_out_valid_filter_5_31,
    hash_out_6_0,
    hash_out_valid_filter_6_0,
    hash_out_6_1,
    hash_out_valid_filter_6_1,
    hash_out_6_2,
    hash_out_valid_filter_6_2,
    hash_out_6_3,
    hash_out_valid_filter_6_3,
    hash_out_6_4,
    hash_out_valid_filter_6_4,
    hash_out_6_5,
    hash_out_valid_filter_6_5,
    hash_out_6_6,
    hash_out_valid_filter_6_6,
    hash_out_6_7,
    hash_out_valid_filter_6_7,
    hash_out_6_8,
    hash_out_valid_filter_6_8,
    hash_out_6_9,
    hash_out_valid_filter_6_9,
    hash_out_6_10,
    hash_out_valid_filter_6_10,
    hash_out_6_11,
    hash_out_valid_filter_6_11,
    hash_out_6_12,
    hash_out_valid_filter_6_12,
    hash_out_6_13,
    hash_out_valid_filter_6_13,
    hash_out_6_14,
    hash_out_valid_filter_6_14,
    hash_out_6_15,
    hash_out_valid_filter_6_15,
    hash_out_6_16,
    hash_out_valid_filter_6_16,
    hash_out_6_17,
    hash_out_valid_filter_6_17,
    hash_out_6_18,
    hash_out_valid_filter_6_18,
    hash_out_6_19,
    hash_out_valid_filter_6_19,
    hash_out_6_20,
    hash_out_valid_filter_6_20,
    hash_out_6_21,
    hash_out_valid_filter_6_21,
    hash_out_6_22,
    hash_out_valid_filter_6_22,
    hash_out_6_23,
    hash_out_valid_filter_6_23,
    hash_out_6_24,
    hash_out_valid_filter_6_24,
    hash_out_6_25,
    hash_out_valid_filter_6_25,
    hash_out_6_26,
    hash_out_valid_filter_6_26,
    hash_out_6_27,
    hash_out_valid_filter_6_27,
    hash_out_6_28,
    hash_out_valid_filter_6_28,
    hash_out_6_29,
    hash_out_valid_filter_6_29,
    hash_out_6_30,
    hash_out_valid_filter_6_30,
    hash_out_6_31,
    hash_out_valid_filter_6_31,
    hash_out_7_0,
    hash_out_valid_filter_7_0,
    hash_out_7_1,
    hash_out_valid_filter_7_1,
    hash_out_7_2,
    hash_out_valid_filter_7_2,
    hash_out_7_3,
    hash_out_valid_filter_7_3,
    hash_out_7_4,
    hash_out_valid_filter_7_4,
    hash_out_7_5,
    hash_out_valid_filter_7_5,
    hash_out_7_6,
    hash_out_valid_filter_7_6,
    hash_out_7_7,
    hash_out_valid_filter_7_7,
    hash_out_7_8,
    hash_out_valid_filter_7_8,
    hash_out_7_9,
    hash_out_valid_filter_7_9,
    hash_out_7_10,
    hash_out_valid_filter_7_10,
    hash_out_7_11,
    hash_out_valid_filter_7_11,
    hash_out_7_12,
    hash_out_valid_filter_7_12,
    hash_out_7_13,
    hash_out_valid_filter_7_13,
    hash_out_7_14,
    hash_out_valid_filter_7_14,
    hash_out_7_15,
    hash_out_valid_filter_7_15,
    hash_out_7_16,
    hash_out_valid_filter_7_16,
    hash_out_7_17,
    hash_out_valid_filter_7_17,
    hash_out_7_18,
    hash_out_valid_filter_7_18,
    hash_out_7_19,
    hash_out_valid_filter_7_19,
    hash_out_7_20,
    hash_out_valid_filter_7_20,
    hash_out_7_21,
    hash_out_valid_filter_7_21,
    hash_out_7_22,
    hash_out_valid_filter_7_22,
    hash_out_7_23,
    hash_out_valid_filter_7_23,
    hash_out_7_24,
    hash_out_valid_filter_7_24,
    hash_out_7_25,
    hash_out_valid_filter_7_25,
    hash_out_7_26,
    hash_out_valid_filter_7_26,
    hash_out_7_27,
    hash_out_valid_filter_7_27,
    hash_out_7_28,
    hash_out_valid_filter_7_28,
    hash_out_7_29,
    hash_out_valid_filter_7_29,
    hash_out_7_30,
    hash_out_valid_filter_7_30,
    hash_out_7_31,
    hash_out_valid_filter_7_31,
    in_data,
    in_valid,
    in_sop,
    in_eop,
    in_empty,
    out_new_pkt
);

input clk;
input rst;
input [255:0] in_data;
input in_valid;
input in_sop;
input in_eop;
input [4:0] in_empty;
output wire [RID_WIDTH-1:0] hash_out_0_0;
output wire hash_out_valid_filter_0_0;
output wire [RID_WIDTH-1:0] hash_out_0_1;
output wire hash_out_valid_filter_0_1;
output wire [RID_WIDTH-1:0] hash_out_0_2;
output wire hash_out_valid_filter_0_2;
output wire [RID_WIDTH-1:0] hash_out_0_3;
output wire hash_out_valid_filter_0_3;
output wire [RID_WIDTH-1:0] hash_out_0_4;
output wire hash_out_valid_filter_0_4;
output wire [RID_WIDTH-1:0] hash_out_0_5;
output wire hash_out_valid_filter_0_5;
output wire [RID_WIDTH-1:0] hash_out_0_6;
output wire hash_out_valid_filter_0_6;
output wire [RID_WIDTH-1:0] hash_out_0_7;
output wire hash_out_valid_filter_0_7;
output wire [RID_WIDTH-1:0] hash_out_0_8;
output wire hash_out_valid_filter_0_8;
output wire [RID_WIDTH-1:0] hash_out_0_9;
output wire hash_out_valid_filter_0_9;
output wire [RID_WIDTH-1:0] hash_out_0_10;
output wire hash_out_valid_filter_0_10;
output wire [RID_WIDTH-1:0] hash_out_0_11;
output wire hash_out_valid_filter_0_11;
output wire [RID_WIDTH-1:0] hash_out_0_12;
output wire hash_out_valid_filter_0_12;
output wire [RID_WIDTH-1:0] hash_out_0_13;
output wire hash_out_valid_filter_0_13;
output wire [RID_WIDTH-1:0] hash_out_0_14;
output wire hash_out_valid_filter_0_14;
output wire [RID_WIDTH-1:0] hash_out_0_15;
output wire hash_out_valid_filter_0_15;
output wire [RID_WIDTH-1:0] hash_out_0_16;
output wire hash_out_valid_filter_0_16;
output wire [RID_WIDTH-1:0] hash_out_0_17;
output wire hash_out_valid_filter_0_17;
output wire [RID_WIDTH-1:0] hash_out_0_18;
output wire hash_out_valid_filter_0_18;
output wire [RID_WIDTH-1:0] hash_out_0_19;
output wire hash_out_valid_filter_0_19;
output wire [RID_WIDTH-1:0] hash_out_0_20;
output wire hash_out_valid_filter_0_20;
output wire [RID_WIDTH-1:0] hash_out_0_21;
output wire hash_out_valid_filter_0_21;
output wire [RID_WIDTH-1:0] hash_out_0_22;
output wire hash_out_valid_filter_0_22;
output wire [RID_WIDTH-1:0] hash_out_0_23;
output wire hash_out_valid_filter_0_23;
output wire [RID_WIDTH-1:0] hash_out_0_24;
output wire hash_out_valid_filter_0_24;
output wire [RID_WIDTH-1:0] hash_out_0_25;
output wire hash_out_valid_filter_0_25;
output wire [RID_WIDTH-1:0] hash_out_0_26;
output wire hash_out_valid_filter_0_26;
output wire [RID_WIDTH-1:0] hash_out_0_27;
output wire hash_out_valid_filter_0_27;
output wire [RID_WIDTH-1:0] hash_out_0_28;
output wire hash_out_valid_filter_0_28;
output wire [RID_WIDTH-1:0] hash_out_0_29;
output wire hash_out_valid_filter_0_29;
output wire [RID_WIDTH-1:0] hash_out_0_30;
output wire hash_out_valid_filter_0_30;
output wire [RID_WIDTH-1:0] hash_out_0_31;
output wire hash_out_valid_filter_0_31;
output wire [RID_WIDTH-1:0] hash_out_1_0;
output wire hash_out_valid_filter_1_0;
output wire [RID_WIDTH-1:0] hash_out_1_1;
output wire hash_out_valid_filter_1_1;
output wire [RID_WIDTH-1:0] hash_out_1_2;
output wire hash_out_valid_filter_1_2;
output wire [RID_WIDTH-1:0] hash_out_1_3;
output wire hash_out_valid_filter_1_3;
output wire [RID_WIDTH-1:0] hash_out_1_4;
output wire hash_out_valid_filter_1_4;
output wire [RID_WIDTH-1:0] hash_out_1_5;
output wire hash_out_valid_filter_1_5;
output wire [RID_WIDTH-1:0] hash_out_1_6;
output wire hash_out_valid_filter_1_6;
output wire [RID_WIDTH-1:0] hash_out_1_7;
output wire hash_out_valid_filter_1_7;
output wire [RID_WIDTH-1:0] hash_out_1_8;
output wire hash_out_valid_filter_1_8;
output wire [RID_WIDTH-1:0] hash_out_1_9;
output wire hash_out_valid_filter_1_9;
output wire [RID_WIDTH-1:0] hash_out_1_10;
output wire hash_out_valid_filter_1_10;
output wire [RID_WIDTH-1:0] hash_out_1_11;
output wire hash_out_valid_filter_1_11;
output wire [RID_WIDTH-1:0] hash_out_1_12;
output wire hash_out_valid_filter_1_12;
output wire [RID_WIDTH-1:0] hash_out_1_13;
output wire hash_out_valid_filter_1_13;
output wire [RID_WIDTH-1:0] hash_out_1_14;
output wire hash_out_valid_filter_1_14;
output wire [RID_WIDTH-1:0] hash_out_1_15;
output wire hash_out_valid_filter_1_15;
output wire [RID_WIDTH-1:0] hash_out_1_16;
output wire hash_out_valid_filter_1_16;
output wire [RID_WIDTH-1:0] hash_out_1_17;
output wire hash_out_valid_filter_1_17;
output wire [RID_WIDTH-1:0] hash_out_1_18;
output wire hash_out_valid_filter_1_18;
output wire [RID_WIDTH-1:0] hash_out_1_19;
output wire hash_out_valid_filter_1_19;
output wire [RID_WIDTH-1:0] hash_out_1_20;
output wire hash_out_valid_filter_1_20;
output wire [RID_WIDTH-1:0] hash_out_1_21;
output wire hash_out_valid_filter_1_21;
output wire [RID_WIDTH-1:0] hash_out_1_22;
output wire hash_out_valid_filter_1_22;
output wire [RID_WIDTH-1:0] hash_out_1_23;
output wire hash_out_valid_filter_1_23;
output wire [RID_WIDTH-1:0] hash_out_1_24;
output wire hash_out_valid_filter_1_24;
output wire [RID_WIDTH-1:0] hash_out_1_25;
output wire hash_out_valid_filter_1_25;
output wire [RID_WIDTH-1:0] hash_out_1_26;
output wire hash_out_valid_filter_1_26;
output wire [RID_WIDTH-1:0] hash_out_1_27;
output wire hash_out_valid_filter_1_27;
output wire [RID_WIDTH-1:0] hash_out_1_28;
output wire hash_out_valid_filter_1_28;
output wire [RID_WIDTH-1:0] hash_out_1_29;
output wire hash_out_valid_filter_1_29;
output wire [RID_WIDTH-1:0] hash_out_1_30;
output wire hash_out_valid_filter_1_30;
output wire [RID_WIDTH-1:0] hash_out_1_31;
output wire hash_out_valid_filter_1_31;
output wire [RID_WIDTH-1:0] hash_out_2_0;
output wire hash_out_valid_filter_2_0;
output wire [RID_WIDTH-1:0] hash_out_2_1;
output wire hash_out_valid_filter_2_1;
output wire [RID_WIDTH-1:0] hash_out_2_2;
output wire hash_out_valid_filter_2_2;
output wire [RID_WIDTH-1:0] hash_out_2_3;
output wire hash_out_valid_filter_2_3;
output wire [RID_WIDTH-1:0] hash_out_2_4;
output wire hash_out_valid_filter_2_4;
output wire [RID_WIDTH-1:0] hash_out_2_5;
output wire hash_out_valid_filter_2_5;
output wire [RID_WIDTH-1:0] hash_out_2_6;
output wire hash_out_valid_filter_2_6;
output wire [RID_WIDTH-1:0] hash_out_2_7;
output wire hash_out_valid_filter_2_7;
output wire [RID_WIDTH-1:0] hash_out_2_8;
output wire hash_out_valid_filter_2_8;
output wire [RID_WIDTH-1:0] hash_out_2_9;
output wire hash_out_valid_filter_2_9;
output wire [RID_WIDTH-1:0] hash_out_2_10;
output wire hash_out_valid_filter_2_10;
output wire [RID_WIDTH-1:0] hash_out_2_11;
output wire hash_out_valid_filter_2_11;
output wire [RID_WIDTH-1:0] hash_out_2_12;
output wire hash_out_valid_filter_2_12;
output wire [RID_WIDTH-1:0] hash_out_2_13;
output wire hash_out_valid_filter_2_13;
output wire [RID_WIDTH-1:0] hash_out_2_14;
output wire hash_out_valid_filter_2_14;
output wire [RID_WIDTH-1:0] hash_out_2_15;
output wire hash_out_valid_filter_2_15;
output wire [RID_WIDTH-1:0] hash_out_2_16;
output wire hash_out_valid_filter_2_16;
output wire [RID_WIDTH-1:0] hash_out_2_17;
output wire hash_out_valid_filter_2_17;
output wire [RID_WIDTH-1:0] hash_out_2_18;
output wire hash_out_valid_filter_2_18;
output wire [RID_WIDTH-1:0] hash_out_2_19;
output wire hash_out_valid_filter_2_19;
output wire [RID_WIDTH-1:0] hash_out_2_20;
output wire hash_out_valid_filter_2_20;
output wire [RID_WIDTH-1:0] hash_out_2_21;
output wire hash_out_valid_filter_2_21;
output wire [RID_WIDTH-1:0] hash_out_2_22;
output wire hash_out_valid_filter_2_22;
output wire [RID_WIDTH-1:0] hash_out_2_23;
output wire hash_out_valid_filter_2_23;
output wire [RID_WIDTH-1:0] hash_out_2_24;
output wire hash_out_valid_filter_2_24;
output wire [RID_WIDTH-1:0] hash_out_2_25;
output wire hash_out_valid_filter_2_25;
output wire [RID_WIDTH-1:0] hash_out_2_26;
output wire hash_out_valid_filter_2_26;
output wire [RID_WIDTH-1:0] hash_out_2_27;
output wire hash_out_valid_filter_2_27;
output wire [RID_WIDTH-1:0] hash_out_2_28;
output wire hash_out_valid_filter_2_28;
output wire [RID_WIDTH-1:0] hash_out_2_29;
output wire hash_out_valid_filter_2_29;
output wire [RID_WIDTH-1:0] hash_out_2_30;
output wire hash_out_valid_filter_2_30;
output wire [RID_WIDTH-1:0] hash_out_2_31;
output wire hash_out_valid_filter_2_31;
output wire [RID_WIDTH-1:0] hash_out_3_0;
output wire hash_out_valid_filter_3_0;
output wire [RID_WIDTH-1:0] hash_out_3_1;
output wire hash_out_valid_filter_3_1;
output wire [RID_WIDTH-1:0] hash_out_3_2;
output wire hash_out_valid_filter_3_2;
output wire [RID_WIDTH-1:0] hash_out_3_3;
output wire hash_out_valid_filter_3_3;
output wire [RID_WIDTH-1:0] hash_out_3_4;
output wire hash_out_valid_filter_3_4;
output wire [RID_WIDTH-1:0] hash_out_3_5;
output wire hash_out_valid_filter_3_5;
output wire [RID_WIDTH-1:0] hash_out_3_6;
output wire hash_out_valid_filter_3_6;
output wire [RID_WIDTH-1:0] hash_out_3_7;
output wire hash_out_valid_filter_3_7;
output wire [RID_WIDTH-1:0] hash_out_3_8;
output wire hash_out_valid_filter_3_8;
output wire [RID_WIDTH-1:0] hash_out_3_9;
output wire hash_out_valid_filter_3_9;
output wire [RID_WIDTH-1:0] hash_out_3_10;
output wire hash_out_valid_filter_3_10;
output wire [RID_WIDTH-1:0] hash_out_3_11;
output wire hash_out_valid_filter_3_11;
output wire [RID_WIDTH-1:0] hash_out_3_12;
output wire hash_out_valid_filter_3_12;
output wire [RID_WIDTH-1:0] hash_out_3_13;
output wire hash_out_valid_filter_3_13;
output wire [RID_WIDTH-1:0] hash_out_3_14;
output wire hash_out_valid_filter_3_14;
output wire [RID_WIDTH-1:0] hash_out_3_15;
output wire hash_out_valid_filter_3_15;
output wire [RID_WIDTH-1:0] hash_out_3_16;
output wire hash_out_valid_filter_3_16;
output wire [RID_WIDTH-1:0] hash_out_3_17;
output wire hash_out_valid_filter_3_17;
output wire [RID_WIDTH-1:0] hash_out_3_18;
output wire hash_out_valid_filter_3_18;
output wire [RID_WIDTH-1:0] hash_out_3_19;
output wire hash_out_valid_filter_3_19;
output wire [RID_WIDTH-1:0] hash_out_3_20;
output wire hash_out_valid_filter_3_20;
output wire [RID_WIDTH-1:0] hash_out_3_21;
output wire hash_out_valid_filter_3_21;
output wire [RID_WIDTH-1:0] hash_out_3_22;
output wire hash_out_valid_filter_3_22;
output wire [RID_WIDTH-1:0] hash_out_3_23;
output wire hash_out_valid_filter_3_23;
output wire [RID_WIDTH-1:0] hash_out_3_24;
output wire hash_out_valid_filter_3_24;
output wire [RID_WIDTH-1:0] hash_out_3_25;
output wire hash_out_valid_filter_3_25;
output wire [RID_WIDTH-1:0] hash_out_3_26;
output wire hash_out_valid_filter_3_26;
output wire [RID_WIDTH-1:0] hash_out_3_27;
output wire hash_out_valid_filter_3_27;
output wire [RID_WIDTH-1:0] hash_out_3_28;
output wire hash_out_valid_filter_3_28;
output wire [RID_WIDTH-1:0] hash_out_3_29;
output wire hash_out_valid_filter_3_29;
output wire [RID_WIDTH-1:0] hash_out_3_30;
output wire hash_out_valid_filter_3_30;
output wire [RID_WIDTH-1:0] hash_out_3_31;
output wire hash_out_valid_filter_3_31;
output wire [RID_WIDTH-1:0] hash_out_4_0;
output wire hash_out_valid_filter_4_0;
output wire [RID_WIDTH-1:0] hash_out_4_1;
output wire hash_out_valid_filter_4_1;
output wire [RID_WIDTH-1:0] hash_out_4_2;
output wire hash_out_valid_filter_4_2;
output wire [RID_WIDTH-1:0] hash_out_4_3;
output wire hash_out_valid_filter_4_3;
output wire [RID_WIDTH-1:0] hash_out_4_4;
output wire hash_out_valid_filter_4_4;
output wire [RID_WIDTH-1:0] hash_out_4_5;
output wire hash_out_valid_filter_4_5;
output wire [RID_WIDTH-1:0] hash_out_4_6;
output wire hash_out_valid_filter_4_6;
output wire [RID_WIDTH-1:0] hash_out_4_7;
output wire hash_out_valid_filter_4_7;
output wire [RID_WIDTH-1:0] hash_out_4_8;
output wire hash_out_valid_filter_4_8;
output wire [RID_WIDTH-1:0] hash_out_4_9;
output wire hash_out_valid_filter_4_9;
output wire [RID_WIDTH-1:0] hash_out_4_10;
output wire hash_out_valid_filter_4_10;
output wire [RID_WIDTH-1:0] hash_out_4_11;
output wire hash_out_valid_filter_4_11;
output wire [RID_WIDTH-1:0] hash_out_4_12;
output wire hash_out_valid_filter_4_12;
output wire [RID_WIDTH-1:0] hash_out_4_13;
output wire hash_out_valid_filter_4_13;
output wire [RID_WIDTH-1:0] hash_out_4_14;
output wire hash_out_valid_filter_4_14;
output wire [RID_WIDTH-1:0] hash_out_4_15;
output wire hash_out_valid_filter_4_15;
output wire [RID_WIDTH-1:0] hash_out_4_16;
output wire hash_out_valid_filter_4_16;
output wire [RID_WIDTH-1:0] hash_out_4_17;
output wire hash_out_valid_filter_4_17;
output wire [RID_WIDTH-1:0] hash_out_4_18;
output wire hash_out_valid_filter_4_18;
output wire [RID_WIDTH-1:0] hash_out_4_19;
output wire hash_out_valid_filter_4_19;
output wire [RID_WIDTH-1:0] hash_out_4_20;
output wire hash_out_valid_filter_4_20;
output wire [RID_WIDTH-1:0] hash_out_4_21;
output wire hash_out_valid_filter_4_21;
output wire [RID_WIDTH-1:0] hash_out_4_22;
output wire hash_out_valid_filter_4_22;
output wire [RID_WIDTH-1:0] hash_out_4_23;
output wire hash_out_valid_filter_4_23;
output wire [RID_WIDTH-1:0] hash_out_4_24;
output wire hash_out_valid_filter_4_24;
output wire [RID_WIDTH-1:0] hash_out_4_25;
output wire hash_out_valid_filter_4_25;
output wire [RID_WIDTH-1:0] hash_out_4_26;
output wire hash_out_valid_filter_4_26;
output wire [RID_WIDTH-1:0] hash_out_4_27;
output wire hash_out_valid_filter_4_27;
output wire [RID_WIDTH-1:0] hash_out_4_28;
output wire hash_out_valid_filter_4_28;
output wire [RID_WIDTH-1:0] hash_out_4_29;
output wire hash_out_valid_filter_4_29;
output wire [RID_WIDTH-1:0] hash_out_4_30;
output wire hash_out_valid_filter_4_30;
output wire [RID_WIDTH-1:0] hash_out_4_31;
output wire hash_out_valid_filter_4_31;
output wire [RID_WIDTH-1:0] hash_out_5_0;
output wire hash_out_valid_filter_5_0;
output wire [RID_WIDTH-1:0] hash_out_5_1;
output wire hash_out_valid_filter_5_1;
output wire [RID_WIDTH-1:0] hash_out_5_2;
output wire hash_out_valid_filter_5_2;
output wire [RID_WIDTH-1:0] hash_out_5_3;
output wire hash_out_valid_filter_5_3;
output wire [RID_WIDTH-1:0] hash_out_5_4;
output wire hash_out_valid_filter_5_4;
output wire [RID_WIDTH-1:0] hash_out_5_5;
output wire hash_out_valid_filter_5_5;
output wire [RID_WIDTH-1:0] hash_out_5_6;
output wire hash_out_valid_filter_5_6;
output wire [RID_WIDTH-1:0] hash_out_5_7;
output wire hash_out_valid_filter_5_7;
output wire [RID_WIDTH-1:0] hash_out_5_8;
output wire hash_out_valid_filter_5_8;
output wire [RID_WIDTH-1:0] hash_out_5_9;
output wire hash_out_valid_filter_5_9;
output wire [RID_WIDTH-1:0] hash_out_5_10;
output wire hash_out_valid_filter_5_10;
output wire [RID_WIDTH-1:0] hash_out_5_11;
output wire hash_out_valid_filter_5_11;
output wire [RID_WIDTH-1:0] hash_out_5_12;
output wire hash_out_valid_filter_5_12;
output wire [RID_WIDTH-1:0] hash_out_5_13;
output wire hash_out_valid_filter_5_13;
output wire [RID_WIDTH-1:0] hash_out_5_14;
output wire hash_out_valid_filter_5_14;
output wire [RID_WIDTH-1:0] hash_out_5_15;
output wire hash_out_valid_filter_5_15;
output wire [RID_WIDTH-1:0] hash_out_5_16;
output wire hash_out_valid_filter_5_16;
output wire [RID_WIDTH-1:0] hash_out_5_17;
output wire hash_out_valid_filter_5_17;
output wire [RID_WIDTH-1:0] hash_out_5_18;
output wire hash_out_valid_filter_5_18;
output wire [RID_WIDTH-1:0] hash_out_5_19;
output wire hash_out_valid_filter_5_19;
output wire [RID_WIDTH-1:0] hash_out_5_20;
output wire hash_out_valid_filter_5_20;
output wire [RID_WIDTH-1:0] hash_out_5_21;
output wire hash_out_valid_filter_5_21;
output wire [RID_WIDTH-1:0] hash_out_5_22;
output wire hash_out_valid_filter_5_22;
output wire [RID_WIDTH-1:0] hash_out_5_23;
output wire hash_out_valid_filter_5_23;
output wire [RID_WIDTH-1:0] hash_out_5_24;
output wire hash_out_valid_filter_5_24;
output wire [RID_WIDTH-1:0] hash_out_5_25;
output wire hash_out_valid_filter_5_25;
output wire [RID_WIDTH-1:0] hash_out_5_26;
output wire hash_out_valid_filter_5_26;
output wire [RID_WIDTH-1:0] hash_out_5_27;
output wire hash_out_valid_filter_5_27;
output wire [RID_WIDTH-1:0] hash_out_5_28;
output wire hash_out_valid_filter_5_28;
output wire [RID_WIDTH-1:0] hash_out_5_29;
output wire hash_out_valid_filter_5_29;
output wire [RID_WIDTH-1:0] hash_out_5_30;
output wire hash_out_valid_filter_5_30;
output wire [RID_WIDTH-1:0] hash_out_5_31;
output wire hash_out_valid_filter_5_31;
output wire [RID_WIDTH-1:0] hash_out_6_0;
output wire hash_out_valid_filter_6_0;
output wire [RID_WIDTH-1:0] hash_out_6_1;
output wire hash_out_valid_filter_6_1;
output wire [RID_WIDTH-1:0] hash_out_6_2;
output wire hash_out_valid_filter_6_2;
output wire [RID_WIDTH-1:0] hash_out_6_3;
output wire hash_out_valid_filter_6_3;
output wire [RID_WIDTH-1:0] hash_out_6_4;
output wire hash_out_valid_filter_6_4;
output wire [RID_WIDTH-1:0] hash_out_6_5;
output wire hash_out_valid_filter_6_5;
output wire [RID_WIDTH-1:0] hash_out_6_6;
output wire hash_out_valid_filter_6_6;
output wire [RID_WIDTH-1:0] hash_out_6_7;
output wire hash_out_valid_filter_6_7;
output wire [RID_WIDTH-1:0] hash_out_6_8;
output wire hash_out_valid_filter_6_8;
output wire [RID_WIDTH-1:0] hash_out_6_9;
output wire hash_out_valid_filter_6_9;
output wire [RID_WIDTH-1:0] hash_out_6_10;
output wire hash_out_valid_filter_6_10;
output wire [RID_WIDTH-1:0] hash_out_6_11;
output wire hash_out_valid_filter_6_11;
output wire [RID_WIDTH-1:0] hash_out_6_12;
output wire hash_out_valid_filter_6_12;
output wire [RID_WIDTH-1:0] hash_out_6_13;
output wire hash_out_valid_filter_6_13;
output wire [RID_WIDTH-1:0] hash_out_6_14;
output wire hash_out_valid_filter_6_14;
output wire [RID_WIDTH-1:0] hash_out_6_15;
output wire hash_out_valid_filter_6_15;
output wire [RID_WIDTH-1:0] hash_out_6_16;
output wire hash_out_valid_filter_6_16;
output wire [RID_WIDTH-1:0] hash_out_6_17;
output wire hash_out_valid_filter_6_17;
output wire [RID_WIDTH-1:0] hash_out_6_18;
output wire hash_out_valid_filter_6_18;
output wire [RID_WIDTH-1:0] hash_out_6_19;
output wire hash_out_valid_filter_6_19;
output wire [RID_WIDTH-1:0] hash_out_6_20;
output wire hash_out_valid_filter_6_20;
output wire [RID_WIDTH-1:0] hash_out_6_21;
output wire hash_out_valid_filter_6_21;
output wire [RID_WIDTH-1:0] hash_out_6_22;
output wire hash_out_valid_filter_6_22;
output wire [RID_WIDTH-1:0] hash_out_6_23;
output wire hash_out_valid_filter_6_23;
output wire [RID_WIDTH-1:0] hash_out_6_24;
output wire hash_out_valid_filter_6_24;
output wire [RID_WIDTH-1:0] hash_out_6_25;
output wire hash_out_valid_filter_6_25;
output wire [RID_WIDTH-1:0] hash_out_6_26;
output wire hash_out_valid_filter_6_26;
output wire [RID_WIDTH-1:0] hash_out_6_27;
output wire hash_out_valid_filter_6_27;
output wire [RID_WIDTH-1:0] hash_out_6_28;
output wire hash_out_valid_filter_6_28;
output wire [RID_WIDTH-1:0] hash_out_6_29;
output wire hash_out_valid_filter_6_29;
output wire [RID_WIDTH-1:0] hash_out_6_30;
output wire hash_out_valid_filter_6_30;
output wire [RID_WIDTH-1:0] hash_out_6_31;
output wire hash_out_valid_filter_6_31;
output wire [RID_WIDTH-1:0] hash_out_7_0;
output wire hash_out_valid_filter_7_0;
output wire [RID_WIDTH-1:0] hash_out_7_1;
output wire hash_out_valid_filter_7_1;
output wire [RID_WIDTH-1:0] hash_out_7_2;
output wire hash_out_valid_filter_7_2;
output wire [RID_WIDTH-1:0] hash_out_7_3;
output wire hash_out_valid_filter_7_3;
output wire [RID_WIDTH-1:0] hash_out_7_4;
output wire hash_out_valid_filter_7_4;
output wire [RID_WIDTH-1:0] hash_out_7_5;
output wire hash_out_valid_filter_7_5;
output wire [RID_WIDTH-1:0] hash_out_7_6;
output wire hash_out_valid_filter_7_6;
output wire [RID_WIDTH-1:0] hash_out_7_7;
output wire hash_out_valid_filter_7_7;
output wire [RID_WIDTH-1:0] hash_out_7_8;
output wire hash_out_valid_filter_7_8;
output wire [RID_WIDTH-1:0] hash_out_7_9;
output wire hash_out_valid_filter_7_9;
output wire [RID_WIDTH-1:0] hash_out_7_10;
output wire hash_out_valid_filter_7_10;
output wire [RID_WIDTH-1:0] hash_out_7_11;
output wire hash_out_valid_filter_7_11;
output wire [RID_WIDTH-1:0] hash_out_7_12;
output wire hash_out_valid_filter_7_12;
output wire [RID_WIDTH-1:0] hash_out_7_13;
output wire hash_out_valid_filter_7_13;
output wire [RID_WIDTH-1:0] hash_out_7_14;
output wire hash_out_valid_filter_7_14;
output wire [RID_WIDTH-1:0] hash_out_7_15;
output wire hash_out_valid_filter_7_15;
output wire [RID_WIDTH-1:0] hash_out_7_16;
output wire hash_out_valid_filter_7_16;
output wire [RID_WIDTH-1:0] hash_out_7_17;
output wire hash_out_valid_filter_7_17;
output wire [RID_WIDTH-1:0] hash_out_7_18;
output wire hash_out_valid_filter_7_18;
output wire [RID_WIDTH-1:0] hash_out_7_19;
output wire hash_out_valid_filter_7_19;
output wire [RID_WIDTH-1:0] hash_out_7_20;
output wire hash_out_valid_filter_7_20;
output wire [RID_WIDTH-1:0] hash_out_7_21;
output wire hash_out_valid_filter_7_21;
output wire [RID_WIDTH-1:0] hash_out_7_22;
output wire hash_out_valid_filter_7_22;
output wire [RID_WIDTH-1:0] hash_out_7_23;
output wire hash_out_valid_filter_7_23;
output wire [RID_WIDTH-1:0] hash_out_7_24;
output wire hash_out_valid_filter_7_24;
output wire [RID_WIDTH-1:0] hash_out_7_25;
output wire hash_out_valid_filter_7_25;
output wire [RID_WIDTH-1:0] hash_out_7_26;
output wire hash_out_valid_filter_7_26;
output wire [RID_WIDTH-1:0] hash_out_7_27;
output wire hash_out_valid_filter_7_27;
output wire [RID_WIDTH-1:0] hash_out_7_28;
output wire hash_out_valid_filter_7_28;
output wire [RID_WIDTH-1:0] hash_out_7_29;
output wire hash_out_valid_filter_7_29;
output wire [RID_WIDTH-1:0] hash_out_7_30;
output wire hash_out_valid_filter_7_30;
output wire [RID_WIDTH-1:0] hash_out_7_31;
output wire hash_out_valid_filter_7_31;
output reg out_new_pkt;

//filter
wire ce;
wire [255:0] filter_out;
wire filter_out_valid;

//hashtable_top
wire hash_out_valid_0_0;
wire hash_out_valid_0_1;
wire hash_out_valid_0_2;
wire hash_out_valid_0_3;
wire hash_out_valid_0_4;
wire hash_out_valid_0_5;
wire hash_out_valid_0_6;
wire hash_out_valid_0_7;
wire hash_out_valid_0_8;
wire hash_out_valid_0_9;
wire hash_out_valid_0_10;
wire hash_out_valid_0_11;
wire hash_out_valid_0_12;
wire hash_out_valid_0_13;
wire hash_out_valid_0_14;
wire hash_out_valid_0_15;
wire hash_out_valid_0_16;
wire hash_out_valid_0_17;
wire hash_out_valid_0_18;
wire hash_out_valid_0_19;
wire hash_out_valid_0_20;
wire hash_out_valid_0_21;
wire hash_out_valid_0_22;
wire hash_out_valid_0_23;
wire hash_out_valid_0_24;
wire hash_out_valid_0_25;
wire hash_out_valid_0_26;
wire hash_out_valid_0_27;
wire hash_out_valid_0_28;
wire hash_out_valid_0_29;
wire hash_out_valid_0_30;
wire hash_out_valid_0_31;
wire hash_out_valid_1_0;
wire hash_out_valid_1_1;
wire hash_out_valid_1_2;
wire hash_out_valid_1_3;
wire hash_out_valid_1_4;
wire hash_out_valid_1_5;
wire hash_out_valid_1_6;
wire hash_out_valid_1_7;
wire hash_out_valid_1_8;
wire hash_out_valid_1_9;
wire hash_out_valid_1_10;
wire hash_out_valid_1_11;
wire hash_out_valid_1_12;
wire hash_out_valid_1_13;
wire hash_out_valid_1_14;
wire hash_out_valid_1_15;
wire hash_out_valid_1_16;
wire hash_out_valid_1_17;
wire hash_out_valid_1_18;
wire hash_out_valid_1_19;
wire hash_out_valid_1_20;
wire hash_out_valid_1_21;
wire hash_out_valid_1_22;
wire hash_out_valid_1_23;
wire hash_out_valid_1_24;
wire hash_out_valid_1_25;
wire hash_out_valid_1_26;
wire hash_out_valid_1_27;
wire hash_out_valid_1_28;
wire hash_out_valid_1_29;
wire hash_out_valid_1_30;
wire hash_out_valid_1_31;
wire hash_out_valid_2_0;
wire hash_out_valid_2_1;
wire hash_out_valid_2_2;
wire hash_out_valid_2_3;
wire hash_out_valid_2_4;
wire hash_out_valid_2_5;
wire hash_out_valid_2_6;
wire hash_out_valid_2_7;
wire hash_out_valid_2_8;
wire hash_out_valid_2_9;
wire hash_out_valid_2_10;
wire hash_out_valid_2_11;
wire hash_out_valid_2_12;
wire hash_out_valid_2_13;
wire hash_out_valid_2_14;
wire hash_out_valid_2_15;
wire hash_out_valid_2_16;
wire hash_out_valid_2_17;
wire hash_out_valid_2_18;
wire hash_out_valid_2_19;
wire hash_out_valid_2_20;
wire hash_out_valid_2_21;
wire hash_out_valid_2_22;
wire hash_out_valid_2_23;
wire hash_out_valid_2_24;
wire hash_out_valid_2_25;
wire hash_out_valid_2_26;
wire hash_out_valid_2_27;
wire hash_out_valid_2_28;
wire hash_out_valid_2_29;
wire hash_out_valid_2_30;
wire hash_out_valid_2_31;
wire hash_out_valid_3_0;
wire hash_out_valid_3_1;
wire hash_out_valid_3_2;
wire hash_out_valid_3_3;
wire hash_out_valid_3_4;
wire hash_out_valid_3_5;
wire hash_out_valid_3_6;
wire hash_out_valid_3_7;
wire hash_out_valid_3_8;
wire hash_out_valid_3_9;
wire hash_out_valid_3_10;
wire hash_out_valid_3_11;
wire hash_out_valid_3_12;
wire hash_out_valid_3_13;
wire hash_out_valid_3_14;
wire hash_out_valid_3_15;
wire hash_out_valid_3_16;
wire hash_out_valid_3_17;
wire hash_out_valid_3_18;
wire hash_out_valid_3_19;
wire hash_out_valid_3_20;
wire hash_out_valid_3_21;
wire hash_out_valid_3_22;
wire hash_out_valid_3_23;
wire hash_out_valid_3_24;
wire hash_out_valid_3_25;
wire hash_out_valid_3_26;
wire hash_out_valid_3_27;
wire hash_out_valid_3_28;
wire hash_out_valid_3_29;
wire hash_out_valid_3_30;
wire hash_out_valid_3_31;
wire hash_out_valid_4_0;
wire hash_out_valid_4_1;
wire hash_out_valid_4_2;
wire hash_out_valid_4_3;
wire hash_out_valid_4_4;
wire hash_out_valid_4_5;
wire hash_out_valid_4_6;
wire hash_out_valid_4_7;
wire hash_out_valid_4_8;
wire hash_out_valid_4_9;
wire hash_out_valid_4_10;
wire hash_out_valid_4_11;
wire hash_out_valid_4_12;
wire hash_out_valid_4_13;
wire hash_out_valid_4_14;
wire hash_out_valid_4_15;
wire hash_out_valid_4_16;
wire hash_out_valid_4_17;
wire hash_out_valid_4_18;
wire hash_out_valid_4_19;
wire hash_out_valid_4_20;
wire hash_out_valid_4_21;
wire hash_out_valid_4_22;
wire hash_out_valid_4_23;
wire hash_out_valid_4_24;
wire hash_out_valid_4_25;
wire hash_out_valid_4_26;
wire hash_out_valid_4_27;
wire hash_out_valid_4_28;
wire hash_out_valid_4_29;
wire hash_out_valid_4_30;
wire hash_out_valid_4_31;
wire hash_out_valid_5_0;
wire hash_out_valid_5_1;
wire hash_out_valid_5_2;
wire hash_out_valid_5_3;
wire hash_out_valid_5_4;
wire hash_out_valid_5_5;
wire hash_out_valid_5_6;
wire hash_out_valid_5_7;
wire hash_out_valid_5_8;
wire hash_out_valid_5_9;
wire hash_out_valid_5_10;
wire hash_out_valid_5_11;
wire hash_out_valid_5_12;
wire hash_out_valid_5_13;
wire hash_out_valid_5_14;
wire hash_out_valid_5_15;
wire hash_out_valid_5_16;
wire hash_out_valid_5_17;
wire hash_out_valid_5_18;
wire hash_out_valid_5_19;
wire hash_out_valid_5_20;
wire hash_out_valid_5_21;
wire hash_out_valid_5_22;
wire hash_out_valid_5_23;
wire hash_out_valid_5_24;
wire hash_out_valid_5_25;
wire hash_out_valid_5_26;
wire hash_out_valid_5_27;
wire hash_out_valid_5_28;
wire hash_out_valid_5_29;
wire hash_out_valid_5_30;
wire hash_out_valid_5_31;
wire hash_out_valid_6_0;
wire hash_out_valid_6_1;
wire hash_out_valid_6_2;
wire hash_out_valid_6_3;
wire hash_out_valid_6_4;
wire hash_out_valid_6_5;
wire hash_out_valid_6_6;
wire hash_out_valid_6_7;
wire hash_out_valid_6_8;
wire hash_out_valid_6_9;
wire hash_out_valid_6_10;
wire hash_out_valid_6_11;
wire hash_out_valid_6_12;
wire hash_out_valid_6_13;
wire hash_out_valid_6_14;
wire hash_out_valid_6_15;
wire hash_out_valid_6_16;
wire hash_out_valid_6_17;
wire hash_out_valid_6_18;
wire hash_out_valid_6_19;
wire hash_out_valid_6_20;
wire hash_out_valid_6_21;
wire hash_out_valid_6_22;
wire hash_out_valid_6_23;
wire hash_out_valid_6_24;
wire hash_out_valid_6_25;
wire hash_out_valid_6_26;
wire hash_out_valid_6_27;
wire hash_out_valid_6_28;
wire hash_out_valid_6_29;
wire hash_out_valid_6_30;
wire hash_out_valid_6_31;
wire hash_out_valid_7_0;
wire hash_out_valid_7_1;
wire hash_out_valid_7_2;
wire hash_out_valid_7_3;
wire hash_out_valid_7_4;
wire hash_out_valid_7_5;
wire hash_out_valid_7_6;
wire hash_out_valid_7_7;
wire hash_out_valid_7_8;
wire hash_out_valid_7_9;
wire hash_out_valid_7_10;
wire hash_out_valid_7_11;
wire hash_out_valid_7_12;
wire hash_out_valid_7_13;
wire hash_out_valid_7_14;
wire hash_out_valid_7_15;
wire hash_out_valid_7_16;
wire hash_out_valid_7_17;
wire hash_out_valid_7_18;
wire hash_out_valid_7_19;
wire hash_out_valid_7_20;
wire hash_out_valid_7_21;
wire hash_out_valid_7_22;
wire hash_out_valid_7_23;
wire hash_out_valid_7_24;
wire hash_out_valid_7_25;
wire hash_out_valid_7_26;
wire hash_out_valid_7_27;
wire hash_out_valid_7_28;
wire hash_out_valid_7_29;
wire hash_out_valid_7_30;
wire hash_out_valid_7_31;
reg [255:0] hash_in;
reg hash_in_valid;

//Other
reg [255:0] din_reg;
reg din_valid_reg;
wire new_pkt;
reg [255:0] filter_out_r1;
reg new_pkt_r1;
reg [255:0] filter_out_r2;
reg new_pkt_r2;
reg [255:0] filter_out_r3;
reg new_pkt_r3;
reg [255:0] filter_out_r4;
reg new_pkt_r4;
reg [255:0] filter_out_r5;
reg new_pkt_r5;
reg [255:0] filter_out_r6;
reg new_pkt_r6;
reg [255:0] filter_out_r7;
reg new_pkt_r7;
reg [255:0] filter_out_r8;
reg new_pkt_r8;
reg [255:0] filter_out_r9;
reg new_pkt_r9;
reg [255:0] filter_out_r10;
reg new_pkt_r10;
reg [255:0] filter_out_r11;
reg new_pkt_r11;
reg [255:0] filter_out_r12;
reg new_pkt_r12;
reg [255:0] filter_out_r13;
reg new_pkt_r13;
reg [255:0] filter_out_r14;
reg new_pkt_r14;
reg [255:0] filter_out_r15;
reg new_pkt_r15;
reg [255:0] filter_out_r16;
reg new_pkt_r16;


`ifdef DUMMY
//No match at all
assign hash_out_valid_filter_0_0 = 0;
assign hash_out_0_0 = 0;
assign hash_out_valid_filter_0_1 = 0;
assign hash_out_0_1 = 0;
assign hash_out_valid_filter_0_2 = 0;
assign hash_out_0_2 = 0;
assign hash_out_valid_filter_0_3 = 0;
assign hash_out_0_3 = 0;
assign hash_out_valid_filter_0_4 = 0;
assign hash_out_0_4 = 0;
assign hash_out_valid_filter_0_5 = 0;
assign hash_out_0_5 = 0;
assign hash_out_valid_filter_0_6 = 0;
assign hash_out_0_6 = 0;
assign hash_out_valid_filter_0_7 = 0;
assign hash_out_0_7 = 0;
assign hash_out_valid_filter_0_8 = 0;
assign hash_out_0_8 = 0;
assign hash_out_valid_filter_0_9 = 0;
assign hash_out_0_9 = 0;
assign hash_out_valid_filter_0_10 = 0;
assign hash_out_0_10 = 0;
assign hash_out_valid_filter_0_11 = 0;
assign hash_out_0_11 = 0;
assign hash_out_valid_filter_0_12 = 0;
assign hash_out_0_12 = 0;
assign hash_out_valid_filter_0_13 = 0;
assign hash_out_0_13 = 0;
assign hash_out_valid_filter_0_14 = 0;
assign hash_out_0_14 = 0;
assign hash_out_valid_filter_0_15 = 0;
assign hash_out_0_15 = 0;
assign hash_out_valid_filter_0_16 = 0;
assign hash_out_0_16 = 0;
assign hash_out_valid_filter_0_17 = 0;
assign hash_out_0_17 = 0;
assign hash_out_valid_filter_0_18 = 0;
assign hash_out_0_18 = 0;
assign hash_out_valid_filter_0_19 = 0;
assign hash_out_0_19 = 0;
assign hash_out_valid_filter_0_20 = 0;
assign hash_out_0_20 = 0;
assign hash_out_valid_filter_0_21 = 0;
assign hash_out_0_21 = 0;
assign hash_out_valid_filter_0_22 = 0;
assign hash_out_0_22 = 0;
assign hash_out_valid_filter_0_23 = 0;
assign hash_out_0_23 = 0;
assign hash_out_valid_filter_0_24 = 0;
assign hash_out_0_24 = 0;
assign hash_out_valid_filter_0_25 = 0;
assign hash_out_0_25 = 0;
assign hash_out_valid_filter_0_26 = 0;
assign hash_out_0_26 = 0;
assign hash_out_valid_filter_0_27 = 0;
assign hash_out_0_27 = 0;
assign hash_out_valid_filter_0_28 = 0;
assign hash_out_0_28 = 0;
assign hash_out_valid_filter_0_29 = 0;
assign hash_out_0_29 = 0;
assign hash_out_valid_filter_0_30 = 0;
assign hash_out_0_30 = 0;
assign hash_out_valid_filter_0_31 = 0;
assign hash_out_0_31 = 0;
assign hash_out_valid_filter_1_0 = 0;
assign hash_out_1_0 = 0;
assign hash_out_valid_filter_1_1 = 0;
assign hash_out_1_1 = 0;
assign hash_out_valid_filter_1_2 = 0;
assign hash_out_1_2 = 0;
assign hash_out_valid_filter_1_3 = 0;
assign hash_out_1_3 = 0;
assign hash_out_valid_filter_1_4 = 0;
assign hash_out_1_4 = 0;
assign hash_out_valid_filter_1_5 = 0;
assign hash_out_1_5 = 0;
assign hash_out_valid_filter_1_6 = 0;
assign hash_out_1_6 = 0;
assign hash_out_valid_filter_1_7 = 0;
assign hash_out_1_7 = 0;
assign hash_out_valid_filter_1_8 = 0;
assign hash_out_1_8 = 0;
assign hash_out_valid_filter_1_9 = 0;
assign hash_out_1_9 = 0;
assign hash_out_valid_filter_1_10 = 0;
assign hash_out_1_10 = 0;
assign hash_out_valid_filter_1_11 = 0;
assign hash_out_1_11 = 0;
assign hash_out_valid_filter_1_12 = 0;
assign hash_out_1_12 = 0;
assign hash_out_valid_filter_1_13 = 0;
assign hash_out_1_13 = 0;
assign hash_out_valid_filter_1_14 = 0;
assign hash_out_1_14 = 0;
assign hash_out_valid_filter_1_15 = 0;
assign hash_out_1_15 = 0;
assign hash_out_valid_filter_1_16 = 0;
assign hash_out_1_16 = 0;
assign hash_out_valid_filter_1_17 = 0;
assign hash_out_1_17 = 0;
assign hash_out_valid_filter_1_18 = 0;
assign hash_out_1_18 = 0;
assign hash_out_valid_filter_1_19 = 0;
assign hash_out_1_19 = 0;
assign hash_out_valid_filter_1_20 = 0;
assign hash_out_1_20 = 0;
assign hash_out_valid_filter_1_21 = 0;
assign hash_out_1_21 = 0;
assign hash_out_valid_filter_1_22 = 0;
assign hash_out_1_22 = 0;
assign hash_out_valid_filter_1_23 = 0;
assign hash_out_1_23 = 0;
assign hash_out_valid_filter_1_24 = 0;
assign hash_out_1_24 = 0;
assign hash_out_valid_filter_1_25 = 0;
assign hash_out_1_25 = 0;
assign hash_out_valid_filter_1_26 = 0;
assign hash_out_1_26 = 0;
assign hash_out_valid_filter_1_27 = 0;
assign hash_out_1_27 = 0;
assign hash_out_valid_filter_1_28 = 0;
assign hash_out_1_28 = 0;
assign hash_out_valid_filter_1_29 = 0;
assign hash_out_1_29 = 0;
assign hash_out_valid_filter_1_30 = 0;
assign hash_out_1_30 = 0;
assign hash_out_valid_filter_1_31 = 0;
assign hash_out_1_31 = 0;
assign hash_out_valid_filter_2_0 = 0;
assign hash_out_2_0 = 0;
assign hash_out_valid_filter_2_1 = 0;
assign hash_out_2_1 = 0;
assign hash_out_valid_filter_2_2 = 0;
assign hash_out_2_2 = 0;
assign hash_out_valid_filter_2_3 = 0;
assign hash_out_2_3 = 0;
assign hash_out_valid_filter_2_4 = 0;
assign hash_out_2_4 = 0;
assign hash_out_valid_filter_2_5 = 0;
assign hash_out_2_5 = 0;
assign hash_out_valid_filter_2_6 = 0;
assign hash_out_2_6 = 0;
assign hash_out_valid_filter_2_7 = 0;
assign hash_out_2_7 = 0;
assign hash_out_valid_filter_2_8 = 0;
assign hash_out_2_8 = 0;
assign hash_out_valid_filter_2_9 = 0;
assign hash_out_2_9 = 0;
assign hash_out_valid_filter_2_10 = 0;
assign hash_out_2_10 = 0;
assign hash_out_valid_filter_2_11 = 0;
assign hash_out_2_11 = 0;
assign hash_out_valid_filter_2_12 = 0;
assign hash_out_2_12 = 0;
assign hash_out_valid_filter_2_13 = 0;
assign hash_out_2_13 = 0;
assign hash_out_valid_filter_2_14 = 0;
assign hash_out_2_14 = 0;
assign hash_out_valid_filter_2_15 = 0;
assign hash_out_2_15 = 0;
assign hash_out_valid_filter_2_16 = 0;
assign hash_out_2_16 = 0;
assign hash_out_valid_filter_2_17 = 0;
assign hash_out_2_17 = 0;
assign hash_out_valid_filter_2_18 = 0;
assign hash_out_2_18 = 0;
assign hash_out_valid_filter_2_19 = 0;
assign hash_out_2_19 = 0;
assign hash_out_valid_filter_2_20 = 0;
assign hash_out_2_20 = 0;
assign hash_out_valid_filter_2_21 = 0;
assign hash_out_2_21 = 0;
assign hash_out_valid_filter_2_22 = 0;
assign hash_out_2_22 = 0;
assign hash_out_valid_filter_2_23 = 0;
assign hash_out_2_23 = 0;
assign hash_out_valid_filter_2_24 = 0;
assign hash_out_2_24 = 0;
assign hash_out_valid_filter_2_25 = 0;
assign hash_out_2_25 = 0;
assign hash_out_valid_filter_2_26 = 0;
assign hash_out_2_26 = 0;
assign hash_out_valid_filter_2_27 = 0;
assign hash_out_2_27 = 0;
assign hash_out_valid_filter_2_28 = 0;
assign hash_out_2_28 = 0;
assign hash_out_valid_filter_2_29 = 0;
assign hash_out_2_29 = 0;
assign hash_out_valid_filter_2_30 = 0;
assign hash_out_2_30 = 0;
assign hash_out_valid_filter_2_31 = 0;
assign hash_out_2_31 = 0;
assign hash_out_valid_filter_3_0 = 0;
assign hash_out_3_0 = 0;
assign hash_out_valid_filter_3_1 = 0;
assign hash_out_3_1 = 0;
assign hash_out_valid_filter_3_2 = 0;
assign hash_out_3_2 = 0;
assign hash_out_valid_filter_3_3 = 0;
assign hash_out_3_3 = 0;
assign hash_out_valid_filter_3_4 = 0;
assign hash_out_3_4 = 0;
assign hash_out_valid_filter_3_5 = 0;
assign hash_out_3_5 = 0;
assign hash_out_valid_filter_3_6 = 0;
assign hash_out_3_6 = 0;
assign hash_out_valid_filter_3_7 = 0;
assign hash_out_3_7 = 0;
assign hash_out_valid_filter_3_8 = 0;
assign hash_out_3_8 = 0;
assign hash_out_valid_filter_3_9 = 0;
assign hash_out_3_9 = 0;
assign hash_out_valid_filter_3_10 = 0;
assign hash_out_3_10 = 0;
assign hash_out_valid_filter_3_11 = 0;
assign hash_out_3_11 = 0;
assign hash_out_valid_filter_3_12 = 0;
assign hash_out_3_12 = 0;
assign hash_out_valid_filter_3_13 = 0;
assign hash_out_3_13 = 0;
assign hash_out_valid_filter_3_14 = 0;
assign hash_out_3_14 = 0;
assign hash_out_valid_filter_3_15 = 0;
assign hash_out_3_15 = 0;
assign hash_out_valid_filter_3_16 = 0;
assign hash_out_3_16 = 0;
assign hash_out_valid_filter_3_17 = 0;
assign hash_out_3_17 = 0;
assign hash_out_valid_filter_3_18 = 0;
assign hash_out_3_18 = 0;
assign hash_out_valid_filter_3_19 = 0;
assign hash_out_3_19 = 0;
assign hash_out_valid_filter_3_20 = 0;
assign hash_out_3_20 = 0;
assign hash_out_valid_filter_3_21 = 0;
assign hash_out_3_21 = 0;
assign hash_out_valid_filter_3_22 = 0;
assign hash_out_3_22 = 0;
assign hash_out_valid_filter_3_23 = 0;
assign hash_out_3_23 = 0;
assign hash_out_valid_filter_3_24 = 0;
assign hash_out_3_24 = 0;
assign hash_out_valid_filter_3_25 = 0;
assign hash_out_3_25 = 0;
assign hash_out_valid_filter_3_26 = 0;
assign hash_out_3_26 = 0;
assign hash_out_valid_filter_3_27 = 0;
assign hash_out_3_27 = 0;
assign hash_out_valid_filter_3_28 = 0;
assign hash_out_3_28 = 0;
assign hash_out_valid_filter_3_29 = 0;
assign hash_out_3_29 = 0;
assign hash_out_valid_filter_3_30 = 0;
assign hash_out_3_30 = 0;
assign hash_out_valid_filter_3_31 = 0;
assign hash_out_3_31 = 0;
assign hash_out_valid_filter_4_0 = 0;
assign hash_out_4_0 = 0;
assign hash_out_valid_filter_4_1 = 0;
assign hash_out_4_1 = 0;
assign hash_out_valid_filter_4_2 = 0;
assign hash_out_4_2 = 0;
assign hash_out_valid_filter_4_3 = 0;
assign hash_out_4_3 = 0;
assign hash_out_valid_filter_4_4 = 0;
assign hash_out_4_4 = 0;
assign hash_out_valid_filter_4_5 = 0;
assign hash_out_4_5 = 0;
assign hash_out_valid_filter_4_6 = 0;
assign hash_out_4_6 = 0;
assign hash_out_valid_filter_4_7 = 0;
assign hash_out_4_7 = 0;
assign hash_out_valid_filter_4_8 = 0;
assign hash_out_4_8 = 0;
assign hash_out_valid_filter_4_9 = 0;
assign hash_out_4_9 = 0;
assign hash_out_valid_filter_4_10 = 0;
assign hash_out_4_10 = 0;
assign hash_out_valid_filter_4_11 = 0;
assign hash_out_4_11 = 0;
assign hash_out_valid_filter_4_12 = 0;
assign hash_out_4_12 = 0;
assign hash_out_valid_filter_4_13 = 0;
assign hash_out_4_13 = 0;
assign hash_out_valid_filter_4_14 = 0;
assign hash_out_4_14 = 0;
assign hash_out_valid_filter_4_15 = 0;
assign hash_out_4_15 = 0;
assign hash_out_valid_filter_4_16 = 0;
assign hash_out_4_16 = 0;
assign hash_out_valid_filter_4_17 = 0;
assign hash_out_4_17 = 0;
assign hash_out_valid_filter_4_18 = 0;
assign hash_out_4_18 = 0;
assign hash_out_valid_filter_4_19 = 0;
assign hash_out_4_19 = 0;
assign hash_out_valid_filter_4_20 = 0;
assign hash_out_4_20 = 0;
assign hash_out_valid_filter_4_21 = 0;
assign hash_out_4_21 = 0;
assign hash_out_valid_filter_4_22 = 0;
assign hash_out_4_22 = 0;
assign hash_out_valid_filter_4_23 = 0;
assign hash_out_4_23 = 0;
assign hash_out_valid_filter_4_24 = 0;
assign hash_out_4_24 = 0;
assign hash_out_valid_filter_4_25 = 0;
assign hash_out_4_25 = 0;
assign hash_out_valid_filter_4_26 = 0;
assign hash_out_4_26 = 0;
assign hash_out_valid_filter_4_27 = 0;
assign hash_out_4_27 = 0;
assign hash_out_valid_filter_4_28 = 0;
assign hash_out_4_28 = 0;
assign hash_out_valid_filter_4_29 = 0;
assign hash_out_4_29 = 0;
assign hash_out_valid_filter_4_30 = 0;
assign hash_out_4_30 = 0;
assign hash_out_valid_filter_4_31 = 0;
assign hash_out_4_31 = 0;
assign hash_out_valid_filter_5_0 = 0;
assign hash_out_5_0 = 0;
assign hash_out_valid_filter_5_1 = 0;
assign hash_out_5_1 = 0;
assign hash_out_valid_filter_5_2 = 0;
assign hash_out_5_2 = 0;
assign hash_out_valid_filter_5_3 = 0;
assign hash_out_5_3 = 0;
assign hash_out_valid_filter_5_4 = 0;
assign hash_out_5_4 = 0;
assign hash_out_valid_filter_5_5 = 0;
assign hash_out_5_5 = 0;
assign hash_out_valid_filter_5_6 = 0;
assign hash_out_5_6 = 0;
assign hash_out_valid_filter_5_7 = 0;
assign hash_out_5_7 = 0;
assign hash_out_valid_filter_5_8 = 0;
assign hash_out_5_8 = 0;
assign hash_out_valid_filter_5_9 = 0;
assign hash_out_5_9 = 0;
assign hash_out_valid_filter_5_10 = 0;
assign hash_out_5_10 = 0;
assign hash_out_valid_filter_5_11 = 0;
assign hash_out_5_11 = 0;
assign hash_out_valid_filter_5_12 = 0;
assign hash_out_5_12 = 0;
assign hash_out_valid_filter_5_13 = 0;
assign hash_out_5_13 = 0;
assign hash_out_valid_filter_5_14 = 0;
assign hash_out_5_14 = 0;
assign hash_out_valid_filter_5_15 = 0;
assign hash_out_5_15 = 0;
assign hash_out_valid_filter_5_16 = 0;
assign hash_out_5_16 = 0;
assign hash_out_valid_filter_5_17 = 0;
assign hash_out_5_17 = 0;
assign hash_out_valid_filter_5_18 = 0;
assign hash_out_5_18 = 0;
assign hash_out_valid_filter_5_19 = 0;
assign hash_out_5_19 = 0;
assign hash_out_valid_filter_5_20 = 0;
assign hash_out_5_20 = 0;
assign hash_out_valid_filter_5_21 = 0;
assign hash_out_5_21 = 0;
assign hash_out_valid_filter_5_22 = 0;
assign hash_out_5_22 = 0;
assign hash_out_valid_filter_5_23 = 0;
assign hash_out_5_23 = 0;
assign hash_out_valid_filter_5_24 = 0;
assign hash_out_5_24 = 0;
assign hash_out_valid_filter_5_25 = 0;
assign hash_out_5_25 = 0;
assign hash_out_valid_filter_5_26 = 0;
assign hash_out_5_26 = 0;
assign hash_out_valid_filter_5_27 = 0;
assign hash_out_5_27 = 0;
assign hash_out_valid_filter_5_28 = 0;
assign hash_out_5_28 = 0;
assign hash_out_valid_filter_5_29 = 0;
assign hash_out_5_29 = 0;
assign hash_out_valid_filter_5_30 = 0;
assign hash_out_5_30 = 0;
assign hash_out_valid_filter_5_31 = 0;
assign hash_out_5_31 = 0;
assign hash_out_valid_filter_6_0 = 0;
assign hash_out_6_0 = 0;
assign hash_out_valid_filter_6_1 = 0;
assign hash_out_6_1 = 0;
assign hash_out_valid_filter_6_2 = 0;
assign hash_out_6_2 = 0;
assign hash_out_valid_filter_6_3 = 0;
assign hash_out_6_3 = 0;
assign hash_out_valid_filter_6_4 = 0;
assign hash_out_6_4 = 0;
assign hash_out_valid_filter_6_5 = 0;
assign hash_out_6_5 = 0;
assign hash_out_valid_filter_6_6 = 0;
assign hash_out_6_6 = 0;
assign hash_out_valid_filter_6_7 = 0;
assign hash_out_6_7 = 0;
assign hash_out_valid_filter_6_8 = 0;
assign hash_out_6_8 = 0;
assign hash_out_valid_filter_6_9 = 0;
assign hash_out_6_9 = 0;
assign hash_out_valid_filter_6_10 = 0;
assign hash_out_6_10 = 0;
assign hash_out_valid_filter_6_11 = 0;
assign hash_out_6_11 = 0;
assign hash_out_valid_filter_6_12 = 0;
assign hash_out_6_12 = 0;
assign hash_out_valid_filter_6_13 = 0;
assign hash_out_6_13 = 0;
assign hash_out_valid_filter_6_14 = 0;
assign hash_out_6_14 = 0;
assign hash_out_valid_filter_6_15 = 0;
assign hash_out_6_15 = 0;
assign hash_out_valid_filter_6_16 = 0;
assign hash_out_6_16 = 0;
assign hash_out_valid_filter_6_17 = 0;
assign hash_out_6_17 = 0;
assign hash_out_valid_filter_6_18 = 0;
assign hash_out_6_18 = 0;
assign hash_out_valid_filter_6_19 = 0;
assign hash_out_6_19 = 0;
assign hash_out_valid_filter_6_20 = 0;
assign hash_out_6_20 = 0;
assign hash_out_valid_filter_6_21 = 0;
assign hash_out_6_21 = 0;
assign hash_out_valid_filter_6_22 = 0;
assign hash_out_6_22 = 0;
assign hash_out_valid_filter_6_23 = 0;
assign hash_out_6_23 = 0;
assign hash_out_valid_filter_6_24 = 0;
assign hash_out_6_24 = 0;
assign hash_out_valid_filter_6_25 = 0;
assign hash_out_6_25 = 0;
assign hash_out_valid_filter_6_26 = 0;
assign hash_out_6_26 = 0;
assign hash_out_valid_filter_6_27 = 0;
assign hash_out_6_27 = 0;
assign hash_out_valid_filter_6_28 = 0;
assign hash_out_6_28 = 0;
assign hash_out_valid_filter_6_29 = 0;
assign hash_out_6_29 = 0;
assign hash_out_valid_filter_6_30 = 0;
assign hash_out_6_30 = 0;
assign hash_out_valid_filter_6_31 = 0;
assign hash_out_6_31 = 0;
assign hash_out_valid_filter_7_0 = 0;
assign hash_out_7_0 = 0;
assign hash_out_valid_filter_7_1 = 0;
assign hash_out_7_1 = 0;
assign hash_out_valid_filter_7_2 = 0;
assign hash_out_7_2 = 0;
assign hash_out_valid_filter_7_3 = 0;
assign hash_out_7_3 = 0;
assign hash_out_valid_filter_7_4 = 0;
assign hash_out_7_4 = 0;
assign hash_out_valid_filter_7_5 = 0;
assign hash_out_7_5 = 0;
assign hash_out_valid_filter_7_6 = 0;
assign hash_out_7_6 = 0;
assign hash_out_valid_filter_7_7 = 0;
assign hash_out_7_7 = 0;
assign hash_out_valid_filter_7_8 = 0;
assign hash_out_7_8 = 0;
assign hash_out_valid_filter_7_9 = 0;
assign hash_out_7_9 = 0;
assign hash_out_valid_filter_7_10 = 0;
assign hash_out_7_10 = 0;
assign hash_out_valid_filter_7_11 = 0;
assign hash_out_7_11 = 0;
assign hash_out_valid_filter_7_12 = 0;
assign hash_out_7_12 = 0;
assign hash_out_valid_filter_7_13 = 0;
assign hash_out_7_13 = 0;
assign hash_out_valid_filter_7_14 = 0;
assign hash_out_7_14 = 0;
assign hash_out_valid_filter_7_15 = 0;
assign hash_out_7_15 = 0;
assign hash_out_valid_filter_7_16 = 0;
assign hash_out_7_16 = 0;
assign hash_out_valid_filter_7_17 = 0;
assign hash_out_7_17 = 0;
assign hash_out_valid_filter_7_18 = 0;
assign hash_out_7_18 = 0;
assign hash_out_valid_filter_7_19 = 0;
assign hash_out_7_19 = 0;
assign hash_out_valid_filter_7_20 = 0;
assign hash_out_7_20 = 0;
assign hash_out_valid_filter_7_21 = 0;
assign hash_out_7_21 = 0;
assign hash_out_valid_filter_7_22 = 0;
assign hash_out_7_22 = 0;
assign hash_out_valid_filter_7_23 = 0;
assign hash_out_7_23 = 0;
assign hash_out_valid_filter_7_24 = 0;
assign hash_out_7_24 = 0;
assign hash_out_valid_filter_7_25 = 0;
assign hash_out_7_25 = 0;
assign hash_out_valid_filter_7_26 = 0;
assign hash_out_7_26 = 0;
assign hash_out_valid_filter_7_27 = 0;
assign hash_out_7_27 = 0;
assign hash_out_valid_filter_7_28 = 0;
assign hash_out_7_28 = 0;
assign hash_out_valid_filter_7_29 = 0;
assign hash_out_7_29 = 0;
assign hash_out_valid_filter_7_30 = 0;
assign hash_out_7_30 = 0;
assign hash_out_valid_filter_7_31 = 0;
assign hash_out_7_31 = 0;

assign new_pkt = in_eop & in_valid;

//Make sure all the flits of the pkts have been checked before moving it. 
always @ (posedge clk) begin
    new_pkt_r1 <= new_pkt;
    new_pkt_r2 <= new_pkt_r1;
    new_pkt_r3 <= new_pkt_r2;
    new_pkt_r4 <= new_pkt_r3;
    new_pkt_r5 <= new_pkt_r4;
    new_pkt_r6 <= new_pkt_r5;
    new_pkt_r7 <= new_pkt_r6;
    new_pkt_r8 <= new_pkt_r7;
    new_pkt_r9 <= new_pkt_r8;
    new_pkt_r10 <= new_pkt_r9;
    new_pkt_r11 <= new_pkt_r10;
    new_pkt_r12 <= new_pkt_r11;
    new_pkt_r13 <= new_pkt_r12;
    new_pkt_r14 <= new_pkt_r13;
    new_pkt_r15 <= new_pkt_r14;
    new_pkt_r16 <= new_pkt_r15;
    out_new_pkt <= new_pkt_r15;
end


`else
//Hashtable signals
assign hash_out_valid_filter_0_0 = hash_out_valid_0_0 & !filter_out_r14[0];
assign hash_out_valid_filter_0_1 = hash_out_valid_0_1 & !filter_out_r14[8];
assign hash_out_valid_filter_0_2 = hash_out_valid_0_2 & !filter_out_r14[16];
assign hash_out_valid_filter_0_3 = hash_out_valid_0_3 & !filter_out_r14[24];
assign hash_out_valid_filter_0_4 = hash_out_valid_0_4 & !filter_out_r14[32];
assign hash_out_valid_filter_0_5 = hash_out_valid_0_5 & !filter_out_r14[40];
assign hash_out_valid_filter_0_6 = hash_out_valid_0_6 & !filter_out_r14[48];
assign hash_out_valid_filter_0_7 = hash_out_valid_0_7 & !filter_out_r14[56];
assign hash_out_valid_filter_0_8 = hash_out_valid_0_8 & !filter_out_r14[64];
assign hash_out_valid_filter_0_9 = hash_out_valid_0_9 & !filter_out_r14[72];
assign hash_out_valid_filter_0_10 = hash_out_valid_0_10 & !filter_out_r14[80];
assign hash_out_valid_filter_0_11 = hash_out_valid_0_11 & !filter_out_r14[88];
assign hash_out_valid_filter_0_12 = hash_out_valid_0_12 & !filter_out_r14[96];
assign hash_out_valid_filter_0_13 = hash_out_valid_0_13 & !filter_out_r14[104];
assign hash_out_valid_filter_0_14 = hash_out_valid_0_14 & !filter_out_r14[112];
assign hash_out_valid_filter_0_15 = hash_out_valid_0_15 & !filter_out_r14[120];
assign hash_out_valid_filter_0_16 = hash_out_valid_0_16 & !filter_out_r14[128];
assign hash_out_valid_filter_0_17 = hash_out_valid_0_17 & !filter_out_r14[136];
assign hash_out_valid_filter_0_18 = hash_out_valid_0_18 & !filter_out_r14[144];
assign hash_out_valid_filter_0_19 = hash_out_valid_0_19 & !filter_out_r14[152];
assign hash_out_valid_filter_0_20 = hash_out_valid_0_20 & !filter_out_r14[160];
assign hash_out_valid_filter_0_21 = hash_out_valid_0_21 & !filter_out_r14[168];
assign hash_out_valid_filter_0_22 = hash_out_valid_0_22 & !filter_out_r14[176];
assign hash_out_valid_filter_0_23 = hash_out_valid_0_23 & !filter_out_r14[184];
assign hash_out_valid_filter_0_24 = hash_out_valid_0_24 & !filter_out_r14[192];
assign hash_out_valid_filter_0_25 = hash_out_valid_0_25 & !filter_out_r14[200];
assign hash_out_valid_filter_0_26 = hash_out_valid_0_26 & !filter_out_r14[208];
assign hash_out_valid_filter_0_27 = hash_out_valid_0_27 & !filter_out_r14[216];
assign hash_out_valid_filter_0_28 = hash_out_valid_0_28 & !filter_out_r14[224];
assign hash_out_valid_filter_0_29 = hash_out_valid_0_29 & !filter_out_r14[232];
assign hash_out_valid_filter_0_30 = hash_out_valid_0_30 & !filter_out_r14[240];
assign hash_out_valid_filter_0_31 = hash_out_valid_0_31 & !filter_out_r14[248];
assign hash_out_valid_filter_1_0 = hash_out_valid_1_0 & !filter_out_r14[1];
assign hash_out_valid_filter_1_1 = hash_out_valid_1_1 & !filter_out_r14[9];
assign hash_out_valid_filter_1_2 = hash_out_valid_1_2 & !filter_out_r14[17];
assign hash_out_valid_filter_1_3 = hash_out_valid_1_3 & !filter_out_r14[25];
assign hash_out_valid_filter_1_4 = hash_out_valid_1_4 & !filter_out_r14[33];
assign hash_out_valid_filter_1_5 = hash_out_valid_1_5 & !filter_out_r14[41];
assign hash_out_valid_filter_1_6 = hash_out_valid_1_6 & !filter_out_r14[49];
assign hash_out_valid_filter_1_7 = hash_out_valid_1_7 & !filter_out_r14[57];
assign hash_out_valid_filter_1_8 = hash_out_valid_1_8 & !filter_out_r14[65];
assign hash_out_valid_filter_1_9 = hash_out_valid_1_9 & !filter_out_r14[73];
assign hash_out_valid_filter_1_10 = hash_out_valid_1_10 & !filter_out_r14[81];
assign hash_out_valid_filter_1_11 = hash_out_valid_1_11 & !filter_out_r14[89];
assign hash_out_valid_filter_1_12 = hash_out_valid_1_12 & !filter_out_r14[97];
assign hash_out_valid_filter_1_13 = hash_out_valid_1_13 & !filter_out_r14[105];
assign hash_out_valid_filter_1_14 = hash_out_valid_1_14 & !filter_out_r14[113];
assign hash_out_valid_filter_1_15 = hash_out_valid_1_15 & !filter_out_r14[121];
assign hash_out_valid_filter_1_16 = hash_out_valid_1_16 & !filter_out_r14[129];
assign hash_out_valid_filter_1_17 = hash_out_valid_1_17 & !filter_out_r14[137];
assign hash_out_valid_filter_1_18 = hash_out_valid_1_18 & !filter_out_r14[145];
assign hash_out_valid_filter_1_19 = hash_out_valid_1_19 & !filter_out_r14[153];
assign hash_out_valid_filter_1_20 = hash_out_valid_1_20 & !filter_out_r14[161];
assign hash_out_valid_filter_1_21 = hash_out_valid_1_21 & !filter_out_r14[169];
assign hash_out_valid_filter_1_22 = hash_out_valid_1_22 & !filter_out_r14[177];
assign hash_out_valid_filter_1_23 = hash_out_valid_1_23 & !filter_out_r14[185];
assign hash_out_valid_filter_1_24 = hash_out_valid_1_24 & !filter_out_r14[193];
assign hash_out_valid_filter_1_25 = hash_out_valid_1_25 & !filter_out_r14[201];
assign hash_out_valid_filter_1_26 = hash_out_valid_1_26 & !filter_out_r14[209];
assign hash_out_valid_filter_1_27 = hash_out_valid_1_27 & !filter_out_r14[217];
assign hash_out_valid_filter_1_28 = hash_out_valid_1_28 & !filter_out_r14[225];
assign hash_out_valid_filter_1_29 = hash_out_valid_1_29 & !filter_out_r14[233];
assign hash_out_valid_filter_1_30 = hash_out_valid_1_30 & !filter_out_r14[241];
assign hash_out_valid_filter_1_31 = hash_out_valid_1_31 & !filter_out_r14[249];
assign hash_out_valid_filter_2_0 = hash_out_valid_2_0 & !filter_out_r14[2];
assign hash_out_valid_filter_2_1 = hash_out_valid_2_1 & !filter_out_r14[10];
assign hash_out_valid_filter_2_2 = hash_out_valid_2_2 & !filter_out_r14[18];
assign hash_out_valid_filter_2_3 = hash_out_valid_2_3 & !filter_out_r14[26];
assign hash_out_valid_filter_2_4 = hash_out_valid_2_4 & !filter_out_r14[34];
assign hash_out_valid_filter_2_5 = hash_out_valid_2_5 & !filter_out_r14[42];
assign hash_out_valid_filter_2_6 = hash_out_valid_2_6 & !filter_out_r14[50];
assign hash_out_valid_filter_2_7 = hash_out_valid_2_7 & !filter_out_r14[58];
assign hash_out_valid_filter_2_8 = hash_out_valid_2_8 & !filter_out_r14[66];
assign hash_out_valid_filter_2_9 = hash_out_valid_2_9 & !filter_out_r14[74];
assign hash_out_valid_filter_2_10 = hash_out_valid_2_10 & !filter_out_r14[82];
assign hash_out_valid_filter_2_11 = hash_out_valid_2_11 & !filter_out_r14[90];
assign hash_out_valid_filter_2_12 = hash_out_valid_2_12 & !filter_out_r14[98];
assign hash_out_valid_filter_2_13 = hash_out_valid_2_13 & !filter_out_r14[106];
assign hash_out_valid_filter_2_14 = hash_out_valid_2_14 & !filter_out_r14[114];
assign hash_out_valid_filter_2_15 = hash_out_valid_2_15 & !filter_out_r14[122];
assign hash_out_valid_filter_2_16 = hash_out_valid_2_16 & !filter_out_r14[130];
assign hash_out_valid_filter_2_17 = hash_out_valid_2_17 & !filter_out_r14[138];
assign hash_out_valid_filter_2_18 = hash_out_valid_2_18 & !filter_out_r14[146];
assign hash_out_valid_filter_2_19 = hash_out_valid_2_19 & !filter_out_r14[154];
assign hash_out_valid_filter_2_20 = hash_out_valid_2_20 & !filter_out_r14[162];
assign hash_out_valid_filter_2_21 = hash_out_valid_2_21 & !filter_out_r14[170];
assign hash_out_valid_filter_2_22 = hash_out_valid_2_22 & !filter_out_r14[178];
assign hash_out_valid_filter_2_23 = hash_out_valid_2_23 & !filter_out_r14[186];
assign hash_out_valid_filter_2_24 = hash_out_valid_2_24 & !filter_out_r14[194];
assign hash_out_valid_filter_2_25 = hash_out_valid_2_25 & !filter_out_r14[202];
assign hash_out_valid_filter_2_26 = hash_out_valid_2_26 & !filter_out_r14[210];
assign hash_out_valid_filter_2_27 = hash_out_valid_2_27 & !filter_out_r14[218];
assign hash_out_valid_filter_2_28 = hash_out_valid_2_28 & !filter_out_r14[226];
assign hash_out_valid_filter_2_29 = hash_out_valid_2_29 & !filter_out_r14[234];
assign hash_out_valid_filter_2_30 = hash_out_valid_2_30 & !filter_out_r14[242];
assign hash_out_valid_filter_2_31 = hash_out_valid_2_31 & !filter_out_r14[250];
assign hash_out_valid_filter_3_0 = hash_out_valid_3_0 & !filter_out_r14[3];
assign hash_out_valid_filter_3_1 = hash_out_valid_3_1 & !filter_out_r14[11];
assign hash_out_valid_filter_3_2 = hash_out_valid_3_2 & !filter_out_r14[19];
assign hash_out_valid_filter_3_3 = hash_out_valid_3_3 & !filter_out_r14[27];
assign hash_out_valid_filter_3_4 = hash_out_valid_3_4 & !filter_out_r14[35];
assign hash_out_valid_filter_3_5 = hash_out_valid_3_5 & !filter_out_r14[43];
assign hash_out_valid_filter_3_6 = hash_out_valid_3_6 & !filter_out_r14[51];
assign hash_out_valid_filter_3_7 = hash_out_valid_3_7 & !filter_out_r14[59];
assign hash_out_valid_filter_3_8 = hash_out_valid_3_8 & !filter_out_r14[67];
assign hash_out_valid_filter_3_9 = hash_out_valid_3_9 & !filter_out_r14[75];
assign hash_out_valid_filter_3_10 = hash_out_valid_3_10 & !filter_out_r14[83];
assign hash_out_valid_filter_3_11 = hash_out_valid_3_11 & !filter_out_r14[91];
assign hash_out_valid_filter_3_12 = hash_out_valid_3_12 & !filter_out_r14[99];
assign hash_out_valid_filter_3_13 = hash_out_valid_3_13 & !filter_out_r14[107];
assign hash_out_valid_filter_3_14 = hash_out_valid_3_14 & !filter_out_r14[115];
assign hash_out_valid_filter_3_15 = hash_out_valid_3_15 & !filter_out_r14[123];
assign hash_out_valid_filter_3_16 = hash_out_valid_3_16 & !filter_out_r14[131];
assign hash_out_valid_filter_3_17 = hash_out_valid_3_17 & !filter_out_r14[139];
assign hash_out_valid_filter_3_18 = hash_out_valid_3_18 & !filter_out_r14[147];
assign hash_out_valid_filter_3_19 = hash_out_valid_3_19 & !filter_out_r14[155];
assign hash_out_valid_filter_3_20 = hash_out_valid_3_20 & !filter_out_r14[163];
assign hash_out_valid_filter_3_21 = hash_out_valid_3_21 & !filter_out_r14[171];
assign hash_out_valid_filter_3_22 = hash_out_valid_3_22 & !filter_out_r14[179];
assign hash_out_valid_filter_3_23 = hash_out_valid_3_23 & !filter_out_r14[187];
assign hash_out_valid_filter_3_24 = hash_out_valid_3_24 & !filter_out_r14[195];
assign hash_out_valid_filter_3_25 = hash_out_valid_3_25 & !filter_out_r14[203];
assign hash_out_valid_filter_3_26 = hash_out_valid_3_26 & !filter_out_r14[211];
assign hash_out_valid_filter_3_27 = hash_out_valid_3_27 & !filter_out_r14[219];
assign hash_out_valid_filter_3_28 = hash_out_valid_3_28 & !filter_out_r14[227];
assign hash_out_valid_filter_3_29 = hash_out_valid_3_29 & !filter_out_r14[235];
assign hash_out_valid_filter_3_30 = hash_out_valid_3_30 & !filter_out_r14[243];
assign hash_out_valid_filter_3_31 = hash_out_valid_3_31 & !filter_out_r14[251];
assign hash_out_valid_filter_4_0 = hash_out_valid_4_0 & !filter_out_r14[4];
assign hash_out_valid_filter_4_1 = hash_out_valid_4_1 & !filter_out_r14[12];
assign hash_out_valid_filter_4_2 = hash_out_valid_4_2 & !filter_out_r14[20];
assign hash_out_valid_filter_4_3 = hash_out_valid_4_3 & !filter_out_r14[28];
assign hash_out_valid_filter_4_4 = hash_out_valid_4_4 & !filter_out_r14[36];
assign hash_out_valid_filter_4_5 = hash_out_valid_4_5 & !filter_out_r14[44];
assign hash_out_valid_filter_4_6 = hash_out_valid_4_6 & !filter_out_r14[52];
assign hash_out_valid_filter_4_7 = hash_out_valid_4_7 & !filter_out_r14[60];
assign hash_out_valid_filter_4_8 = hash_out_valid_4_8 & !filter_out_r14[68];
assign hash_out_valid_filter_4_9 = hash_out_valid_4_9 & !filter_out_r14[76];
assign hash_out_valid_filter_4_10 = hash_out_valid_4_10 & !filter_out_r14[84];
assign hash_out_valid_filter_4_11 = hash_out_valid_4_11 & !filter_out_r14[92];
assign hash_out_valid_filter_4_12 = hash_out_valid_4_12 & !filter_out_r14[100];
assign hash_out_valid_filter_4_13 = hash_out_valid_4_13 & !filter_out_r14[108];
assign hash_out_valid_filter_4_14 = hash_out_valid_4_14 & !filter_out_r14[116];
assign hash_out_valid_filter_4_15 = hash_out_valid_4_15 & !filter_out_r14[124];
assign hash_out_valid_filter_4_16 = hash_out_valid_4_16 & !filter_out_r14[132];
assign hash_out_valid_filter_4_17 = hash_out_valid_4_17 & !filter_out_r14[140];
assign hash_out_valid_filter_4_18 = hash_out_valid_4_18 & !filter_out_r14[148];
assign hash_out_valid_filter_4_19 = hash_out_valid_4_19 & !filter_out_r14[156];
assign hash_out_valid_filter_4_20 = hash_out_valid_4_20 & !filter_out_r14[164];
assign hash_out_valid_filter_4_21 = hash_out_valid_4_21 & !filter_out_r14[172];
assign hash_out_valid_filter_4_22 = hash_out_valid_4_22 & !filter_out_r14[180];
assign hash_out_valid_filter_4_23 = hash_out_valid_4_23 & !filter_out_r14[188];
assign hash_out_valid_filter_4_24 = hash_out_valid_4_24 & !filter_out_r14[196];
assign hash_out_valid_filter_4_25 = hash_out_valid_4_25 & !filter_out_r14[204];
assign hash_out_valid_filter_4_26 = hash_out_valid_4_26 & !filter_out_r14[212];
assign hash_out_valid_filter_4_27 = hash_out_valid_4_27 & !filter_out_r14[220];
assign hash_out_valid_filter_4_28 = hash_out_valid_4_28 & !filter_out_r14[228];
assign hash_out_valid_filter_4_29 = hash_out_valid_4_29 & !filter_out_r14[236];
assign hash_out_valid_filter_4_30 = hash_out_valid_4_30 & !filter_out_r14[244];
assign hash_out_valid_filter_4_31 = hash_out_valid_4_31 & !filter_out_r14[252];
assign hash_out_valid_filter_5_0 = hash_out_valid_5_0 & !filter_out_r14[5];
assign hash_out_valid_filter_5_1 = hash_out_valid_5_1 & !filter_out_r14[13];
assign hash_out_valid_filter_5_2 = hash_out_valid_5_2 & !filter_out_r14[21];
assign hash_out_valid_filter_5_3 = hash_out_valid_5_3 & !filter_out_r14[29];
assign hash_out_valid_filter_5_4 = hash_out_valid_5_4 & !filter_out_r14[37];
assign hash_out_valid_filter_5_5 = hash_out_valid_5_5 & !filter_out_r14[45];
assign hash_out_valid_filter_5_6 = hash_out_valid_5_6 & !filter_out_r14[53];
assign hash_out_valid_filter_5_7 = hash_out_valid_5_7 & !filter_out_r14[61];
assign hash_out_valid_filter_5_8 = hash_out_valid_5_8 & !filter_out_r14[69];
assign hash_out_valid_filter_5_9 = hash_out_valid_5_9 & !filter_out_r14[77];
assign hash_out_valid_filter_5_10 = hash_out_valid_5_10 & !filter_out_r14[85];
assign hash_out_valid_filter_5_11 = hash_out_valid_5_11 & !filter_out_r14[93];
assign hash_out_valid_filter_5_12 = hash_out_valid_5_12 & !filter_out_r14[101];
assign hash_out_valid_filter_5_13 = hash_out_valid_5_13 & !filter_out_r14[109];
assign hash_out_valid_filter_5_14 = hash_out_valid_5_14 & !filter_out_r14[117];
assign hash_out_valid_filter_5_15 = hash_out_valid_5_15 & !filter_out_r14[125];
assign hash_out_valid_filter_5_16 = hash_out_valid_5_16 & !filter_out_r14[133];
assign hash_out_valid_filter_5_17 = hash_out_valid_5_17 & !filter_out_r14[141];
assign hash_out_valid_filter_5_18 = hash_out_valid_5_18 & !filter_out_r14[149];
assign hash_out_valid_filter_5_19 = hash_out_valid_5_19 & !filter_out_r14[157];
assign hash_out_valid_filter_5_20 = hash_out_valid_5_20 & !filter_out_r14[165];
assign hash_out_valid_filter_5_21 = hash_out_valid_5_21 & !filter_out_r14[173];
assign hash_out_valid_filter_5_22 = hash_out_valid_5_22 & !filter_out_r14[181];
assign hash_out_valid_filter_5_23 = hash_out_valid_5_23 & !filter_out_r14[189];
assign hash_out_valid_filter_5_24 = hash_out_valid_5_24 & !filter_out_r14[197];
assign hash_out_valid_filter_5_25 = hash_out_valid_5_25 & !filter_out_r14[205];
assign hash_out_valid_filter_5_26 = hash_out_valid_5_26 & !filter_out_r14[213];
assign hash_out_valid_filter_5_27 = hash_out_valid_5_27 & !filter_out_r14[221];
assign hash_out_valid_filter_5_28 = hash_out_valid_5_28 & !filter_out_r14[229];
assign hash_out_valid_filter_5_29 = hash_out_valid_5_29 & !filter_out_r14[237];
assign hash_out_valid_filter_5_30 = hash_out_valid_5_30 & !filter_out_r14[245];
assign hash_out_valid_filter_5_31 = hash_out_valid_5_31 & !filter_out_r14[253];
assign hash_out_valid_filter_6_0 = hash_out_valid_6_0 & !filter_out_r14[6];
assign hash_out_valid_filter_6_1 = hash_out_valid_6_1 & !filter_out_r14[14];
assign hash_out_valid_filter_6_2 = hash_out_valid_6_2 & !filter_out_r14[22];
assign hash_out_valid_filter_6_3 = hash_out_valid_6_3 & !filter_out_r14[30];
assign hash_out_valid_filter_6_4 = hash_out_valid_6_4 & !filter_out_r14[38];
assign hash_out_valid_filter_6_5 = hash_out_valid_6_5 & !filter_out_r14[46];
assign hash_out_valid_filter_6_6 = hash_out_valid_6_6 & !filter_out_r14[54];
assign hash_out_valid_filter_6_7 = hash_out_valid_6_7 & !filter_out_r14[62];
assign hash_out_valid_filter_6_8 = hash_out_valid_6_8 & !filter_out_r14[70];
assign hash_out_valid_filter_6_9 = hash_out_valid_6_9 & !filter_out_r14[78];
assign hash_out_valid_filter_6_10 = hash_out_valid_6_10 & !filter_out_r14[86];
assign hash_out_valid_filter_6_11 = hash_out_valid_6_11 & !filter_out_r14[94];
assign hash_out_valid_filter_6_12 = hash_out_valid_6_12 & !filter_out_r14[102];
assign hash_out_valid_filter_6_13 = hash_out_valid_6_13 & !filter_out_r14[110];
assign hash_out_valid_filter_6_14 = hash_out_valid_6_14 & !filter_out_r14[118];
assign hash_out_valid_filter_6_15 = hash_out_valid_6_15 & !filter_out_r14[126];
assign hash_out_valid_filter_6_16 = hash_out_valid_6_16 & !filter_out_r14[134];
assign hash_out_valid_filter_6_17 = hash_out_valid_6_17 & !filter_out_r14[142];
assign hash_out_valid_filter_6_18 = hash_out_valid_6_18 & !filter_out_r14[150];
assign hash_out_valid_filter_6_19 = hash_out_valid_6_19 & !filter_out_r14[158];
assign hash_out_valid_filter_6_20 = hash_out_valid_6_20 & !filter_out_r14[166];
assign hash_out_valid_filter_6_21 = hash_out_valid_6_21 & !filter_out_r14[174];
assign hash_out_valid_filter_6_22 = hash_out_valid_6_22 & !filter_out_r14[182];
assign hash_out_valid_filter_6_23 = hash_out_valid_6_23 & !filter_out_r14[190];
assign hash_out_valid_filter_6_24 = hash_out_valid_6_24 & !filter_out_r14[198];
assign hash_out_valid_filter_6_25 = hash_out_valid_6_25 & !filter_out_r14[206];
assign hash_out_valid_filter_6_26 = hash_out_valid_6_26 & !filter_out_r14[214];
assign hash_out_valid_filter_6_27 = hash_out_valid_6_27 & !filter_out_r14[222];
assign hash_out_valid_filter_6_28 = hash_out_valid_6_28 & !filter_out_r14[230];
assign hash_out_valid_filter_6_29 = hash_out_valid_6_29 & !filter_out_r14[238];
assign hash_out_valid_filter_6_30 = hash_out_valid_6_30 & !filter_out_r14[246];
assign hash_out_valid_filter_6_31 = hash_out_valid_6_31 & !filter_out_r14[254];
assign hash_out_valid_filter_7_0 = hash_out_valid_7_0 & !filter_out_r14[7];
assign hash_out_valid_filter_7_1 = hash_out_valid_7_1 & !filter_out_r14[15];
assign hash_out_valid_filter_7_2 = hash_out_valid_7_2 & !filter_out_r14[23];
assign hash_out_valid_filter_7_3 = hash_out_valid_7_3 & !filter_out_r14[31];
assign hash_out_valid_filter_7_4 = hash_out_valid_7_4 & !filter_out_r14[39];
assign hash_out_valid_filter_7_5 = hash_out_valid_7_5 & !filter_out_r14[47];
assign hash_out_valid_filter_7_6 = hash_out_valid_7_6 & !filter_out_r14[55];
assign hash_out_valid_filter_7_7 = hash_out_valid_7_7 & !filter_out_r14[63];
assign hash_out_valid_filter_7_8 = hash_out_valid_7_8 & !filter_out_r14[71];
assign hash_out_valid_filter_7_9 = hash_out_valid_7_9 & !filter_out_r14[79];
assign hash_out_valid_filter_7_10 = hash_out_valid_7_10 & !filter_out_r14[87];
assign hash_out_valid_filter_7_11 = hash_out_valid_7_11 & !filter_out_r14[95];
assign hash_out_valid_filter_7_12 = hash_out_valid_7_12 & !filter_out_r14[103];
assign hash_out_valid_filter_7_13 = hash_out_valid_7_13 & !filter_out_r14[111];
assign hash_out_valid_filter_7_14 = hash_out_valid_7_14 & !filter_out_r14[119];
assign hash_out_valid_filter_7_15 = hash_out_valid_7_15 & !filter_out_r14[127];
assign hash_out_valid_filter_7_16 = hash_out_valid_7_16 & !filter_out_r14[135];
assign hash_out_valid_filter_7_17 = hash_out_valid_7_17 & !filter_out_r14[143];
assign hash_out_valid_filter_7_18 = hash_out_valid_7_18 & !filter_out_r14[151];
assign hash_out_valid_filter_7_19 = hash_out_valid_7_19 & !filter_out_r14[159];
assign hash_out_valid_filter_7_20 = hash_out_valid_7_20 & !filter_out_r14[167];
assign hash_out_valid_filter_7_21 = hash_out_valid_7_21 & !filter_out_r14[175];
assign hash_out_valid_filter_7_22 = hash_out_valid_7_22 & !filter_out_r14[183];
assign hash_out_valid_filter_7_23 = hash_out_valid_7_23 & !filter_out_r14[191];
assign hash_out_valid_filter_7_24 = hash_out_valid_7_24 & !filter_out_r14[199];
assign hash_out_valid_filter_7_25 = hash_out_valid_7_25 & !filter_out_r14[207];
assign hash_out_valid_filter_7_26 = hash_out_valid_7_26 & !filter_out_r14[215];
assign hash_out_valid_filter_7_27 = hash_out_valid_7_27 & !filter_out_r14[223];
assign hash_out_valid_filter_7_28 = hash_out_valid_7_28 & !filter_out_r14[231];
assign hash_out_valid_filter_7_29 = hash_out_valid_7_29 & !filter_out_r14[239];
assign hash_out_valid_filter_7_30 = hash_out_valid_7_30 & !filter_out_r14[247];
assign hash_out_valid_filter_7_31 = hash_out_valid_7_31 & !filter_out_r14[255];

assign new_pkt = in_eop & in_valid;

//Make sure all the flits of the pkts have been checked before moving it. 
always @ (posedge clk) begin
    //if(rst) begin
    //    out_new_pkt <= 0;
    //    new_pkt_r1 <= 0;
    //    new_pkt_r2 <= 0;
    //    new_pkt_r3 <= 0;
    //    new_pkt_r4 <= 0;
    //    new_pkt_r5 <= 0;
    //    new_pkt_r6 <= 0;
    //    new_pkt_r7 <= 0;
    //    new_pkt_r8 <= 0;
    //    new_pkt_r9 <= 0;
    //    new_pkt_r10 <= 0;
    //    new_pkt_r11 <= 0;
    //    new_pkt_r12 <= 0;
    //    new_pkt_r13 <= 0;
    //    new_pkt_r14 <= 0;
    //    new_pkt_r15 <= 0;
    //    new_pkt_r16 <= 0;
    //end else begin
        new_pkt_r1 <= new_pkt;
        new_pkt_r2 <= new_pkt_r1;
        new_pkt_r3 <= new_pkt_r2;
        new_pkt_r4 <= new_pkt_r3;
        new_pkt_r5 <= new_pkt_r4;
        new_pkt_r6 <= new_pkt_r5;
        new_pkt_r7 <= new_pkt_r6;
        new_pkt_r8 <= new_pkt_r7;
        new_pkt_r9 <= new_pkt_r8;
        new_pkt_r10 <= new_pkt_r9;
        new_pkt_r11 <= new_pkt_r10;
        new_pkt_r12 <= new_pkt_r11;
        new_pkt_r13 <= new_pkt_r12;
        new_pkt_r14 <= new_pkt_r13;
        new_pkt_r15 <= new_pkt_r14;
        new_pkt_r16 <= new_pkt_r15;
        out_new_pkt <= new_pkt_r15;
    //end
end

//consistent with the filter 
always @ (posedge clk) begin
    hash_in <= in_data;
    hash_in_valid <= in_valid;
end


//Comb of filter and hashtable
always @ (posedge clk) begin
    //if(rst) begin
    //    filter_out_r1 <= {256{1'b1}};
    //    filter_out_r2 <= {256{1'b1}};
    //    filter_out_r3 <= {256{1'b1}};
    //    filter_out_r4 <= {256{1'b1}};
    //    filter_out_r5 <= {256{1'b1}};
    //    filter_out_r6 <= {256{1'b1}};
    //    filter_out_r7 <= {256{1'b1}};
    //    filter_out_r8 <= {256{1'b1}};
    //    filter_out_r9 <= {256{1'b1}};
    //    filter_out_r10 <= {256{1'b1}};
    //    filter_out_r11 <= {256{1'b1}};
    //    filter_out_r12 <= {256{1'b1}};
    //    filter_out_r13 <= {256{1'b1}};
    //    filter_out_r14 <= {256{1'b1}};
    //    filter_out_r15 <= {256{1'b1}};
    //end else begin
        if(filter_out_valid) begin
            filter_out_r1 <= filter_out;
        end else begin
            filter_out_r1 <= {256{1'b1}};
        end
        filter_out_r2 <= filter_out_r1;
        filter_out_r3 <= filter_out_r2;
        filter_out_r4 <= filter_out_r3;
        filter_out_r5 <= filter_out_r4;
        filter_out_r6 <= filter_out_r5;
        filter_out_r7 <= filter_out_r6;
        filter_out_r8 <= filter_out_r7;
        filter_out_r9 <= filter_out_r8;
        filter_out_r10 <= filter_out_r9;
        filter_out_r11 <= filter_out_r10;
        filter_out_r12 <= filter_out_r11;
        filter_out_r13 <= filter_out_r12;
        filter_out_r14 <= filter_out_r13;
    //end
end


//Instantiation
first_filter filter_inst(
    .clk(clk),
    .rst(rst),
	.in_data    (in_data),
    .in_valid   (in_valid),
    .in_sop     (in_sop),
    .in_eop     (in_eop),
    .in_empty   (in_empty),
    .out_data   (filter_out),
    .out_valid  (filter_out_valid)
);

hashtable_top hashtable_top_inst (
	.clk (clk),
	.dout_0_0 (hash_out_0_0),
    .dout_valid_0_0 (hash_out_valid_0_0),
	.dout_0_1 (hash_out_0_1),
    .dout_valid_0_1 (hash_out_valid_0_1),
	.dout_0_2 (hash_out_0_2),
    .dout_valid_0_2 (hash_out_valid_0_2),
	.dout_0_3 (hash_out_0_3),
    .dout_valid_0_3 (hash_out_valid_0_3),
	.dout_0_4 (hash_out_0_4),
    .dout_valid_0_4 (hash_out_valid_0_4),
	.dout_0_5 (hash_out_0_5),
    .dout_valid_0_5 (hash_out_valid_0_5),
	.dout_0_6 (hash_out_0_6),
    .dout_valid_0_6 (hash_out_valid_0_6),
	.dout_0_7 (hash_out_0_7),
    .dout_valid_0_7 (hash_out_valid_0_7),
	.dout_0_8 (hash_out_0_8),
    .dout_valid_0_8 (hash_out_valid_0_8),
	.dout_0_9 (hash_out_0_9),
    .dout_valid_0_9 (hash_out_valid_0_9),
	.dout_0_10 (hash_out_0_10),
    .dout_valid_0_10 (hash_out_valid_0_10),
	.dout_0_11 (hash_out_0_11),
    .dout_valid_0_11 (hash_out_valid_0_11),
	.dout_0_12 (hash_out_0_12),
    .dout_valid_0_12 (hash_out_valid_0_12),
	.dout_0_13 (hash_out_0_13),
    .dout_valid_0_13 (hash_out_valid_0_13),
	.dout_0_14 (hash_out_0_14),
    .dout_valid_0_14 (hash_out_valid_0_14),
	.dout_0_15 (hash_out_0_15),
    .dout_valid_0_15 (hash_out_valid_0_15),
	.dout_0_16 (hash_out_0_16),
    .dout_valid_0_16 (hash_out_valid_0_16),
	.dout_0_17 (hash_out_0_17),
    .dout_valid_0_17 (hash_out_valid_0_17),
	.dout_0_18 (hash_out_0_18),
    .dout_valid_0_18 (hash_out_valid_0_18),
	.dout_0_19 (hash_out_0_19),
    .dout_valid_0_19 (hash_out_valid_0_19),
	.dout_0_20 (hash_out_0_20),
    .dout_valid_0_20 (hash_out_valid_0_20),
	.dout_0_21 (hash_out_0_21),
    .dout_valid_0_21 (hash_out_valid_0_21),
	.dout_0_22 (hash_out_0_22),
    .dout_valid_0_22 (hash_out_valid_0_22),
	.dout_0_23 (hash_out_0_23),
    .dout_valid_0_23 (hash_out_valid_0_23),
	.dout_0_24 (hash_out_0_24),
    .dout_valid_0_24 (hash_out_valid_0_24),
	.dout_0_25 (hash_out_0_25),
    .dout_valid_0_25 (hash_out_valid_0_25),
	.dout_0_26 (hash_out_0_26),
    .dout_valid_0_26 (hash_out_valid_0_26),
	.dout_0_27 (hash_out_0_27),
    .dout_valid_0_27 (hash_out_valid_0_27),
	.dout_0_28 (hash_out_0_28),
    .dout_valid_0_28 (hash_out_valid_0_28),
	.dout_0_29 (hash_out_0_29),
    .dout_valid_0_29 (hash_out_valid_0_29),
	.dout_0_30 (hash_out_0_30),
    .dout_valid_0_30 (hash_out_valid_0_30),
	.dout_0_31 (hash_out_0_31),
    .dout_valid_0_31 (hash_out_valid_0_31),
	.dout_1_0 (hash_out_1_0),
    .dout_valid_1_0 (hash_out_valid_1_0),
	.dout_1_1 (hash_out_1_1),
    .dout_valid_1_1 (hash_out_valid_1_1),
	.dout_1_2 (hash_out_1_2),
    .dout_valid_1_2 (hash_out_valid_1_2),
	.dout_1_3 (hash_out_1_3),
    .dout_valid_1_3 (hash_out_valid_1_3),
	.dout_1_4 (hash_out_1_4),
    .dout_valid_1_4 (hash_out_valid_1_4),
	.dout_1_5 (hash_out_1_5),
    .dout_valid_1_5 (hash_out_valid_1_5),
	.dout_1_6 (hash_out_1_6),
    .dout_valid_1_6 (hash_out_valid_1_6),
	.dout_1_7 (hash_out_1_7),
    .dout_valid_1_7 (hash_out_valid_1_7),
	.dout_1_8 (hash_out_1_8),
    .dout_valid_1_8 (hash_out_valid_1_8),
	.dout_1_9 (hash_out_1_9),
    .dout_valid_1_9 (hash_out_valid_1_9),
	.dout_1_10 (hash_out_1_10),
    .dout_valid_1_10 (hash_out_valid_1_10),
	.dout_1_11 (hash_out_1_11),
    .dout_valid_1_11 (hash_out_valid_1_11),
	.dout_1_12 (hash_out_1_12),
    .dout_valid_1_12 (hash_out_valid_1_12),
	.dout_1_13 (hash_out_1_13),
    .dout_valid_1_13 (hash_out_valid_1_13),
	.dout_1_14 (hash_out_1_14),
    .dout_valid_1_14 (hash_out_valid_1_14),
	.dout_1_15 (hash_out_1_15),
    .dout_valid_1_15 (hash_out_valid_1_15),
	.dout_1_16 (hash_out_1_16),
    .dout_valid_1_16 (hash_out_valid_1_16),
	.dout_1_17 (hash_out_1_17),
    .dout_valid_1_17 (hash_out_valid_1_17),
	.dout_1_18 (hash_out_1_18),
    .dout_valid_1_18 (hash_out_valid_1_18),
	.dout_1_19 (hash_out_1_19),
    .dout_valid_1_19 (hash_out_valid_1_19),
	.dout_1_20 (hash_out_1_20),
    .dout_valid_1_20 (hash_out_valid_1_20),
	.dout_1_21 (hash_out_1_21),
    .dout_valid_1_21 (hash_out_valid_1_21),
	.dout_1_22 (hash_out_1_22),
    .dout_valid_1_22 (hash_out_valid_1_22),
	.dout_1_23 (hash_out_1_23),
    .dout_valid_1_23 (hash_out_valid_1_23),
	.dout_1_24 (hash_out_1_24),
    .dout_valid_1_24 (hash_out_valid_1_24),
	.dout_1_25 (hash_out_1_25),
    .dout_valid_1_25 (hash_out_valid_1_25),
	.dout_1_26 (hash_out_1_26),
    .dout_valid_1_26 (hash_out_valid_1_26),
	.dout_1_27 (hash_out_1_27),
    .dout_valid_1_27 (hash_out_valid_1_27),
	.dout_1_28 (hash_out_1_28),
    .dout_valid_1_28 (hash_out_valid_1_28),
	.dout_1_29 (hash_out_1_29),
    .dout_valid_1_29 (hash_out_valid_1_29),
	.dout_1_30 (hash_out_1_30),
    .dout_valid_1_30 (hash_out_valid_1_30),
	.dout_1_31 (hash_out_1_31),
    .dout_valid_1_31 (hash_out_valid_1_31),
	.dout_2_0 (hash_out_2_0),
    .dout_valid_2_0 (hash_out_valid_2_0),
	.dout_2_1 (hash_out_2_1),
    .dout_valid_2_1 (hash_out_valid_2_1),
	.dout_2_2 (hash_out_2_2),
    .dout_valid_2_2 (hash_out_valid_2_2),
	.dout_2_3 (hash_out_2_3),
    .dout_valid_2_3 (hash_out_valid_2_3),
	.dout_2_4 (hash_out_2_4),
    .dout_valid_2_4 (hash_out_valid_2_4),
	.dout_2_5 (hash_out_2_5),
    .dout_valid_2_5 (hash_out_valid_2_5),
	.dout_2_6 (hash_out_2_6),
    .dout_valid_2_6 (hash_out_valid_2_6),
	.dout_2_7 (hash_out_2_7),
    .dout_valid_2_7 (hash_out_valid_2_7),
	.dout_2_8 (hash_out_2_8),
    .dout_valid_2_8 (hash_out_valid_2_8),
	.dout_2_9 (hash_out_2_9),
    .dout_valid_2_9 (hash_out_valid_2_9),
	.dout_2_10 (hash_out_2_10),
    .dout_valid_2_10 (hash_out_valid_2_10),
	.dout_2_11 (hash_out_2_11),
    .dout_valid_2_11 (hash_out_valid_2_11),
	.dout_2_12 (hash_out_2_12),
    .dout_valid_2_12 (hash_out_valid_2_12),
	.dout_2_13 (hash_out_2_13),
    .dout_valid_2_13 (hash_out_valid_2_13),
	.dout_2_14 (hash_out_2_14),
    .dout_valid_2_14 (hash_out_valid_2_14),
	.dout_2_15 (hash_out_2_15),
    .dout_valid_2_15 (hash_out_valid_2_15),
	.dout_2_16 (hash_out_2_16),
    .dout_valid_2_16 (hash_out_valid_2_16),
	.dout_2_17 (hash_out_2_17),
    .dout_valid_2_17 (hash_out_valid_2_17),
	.dout_2_18 (hash_out_2_18),
    .dout_valid_2_18 (hash_out_valid_2_18),
	.dout_2_19 (hash_out_2_19),
    .dout_valid_2_19 (hash_out_valid_2_19),
	.dout_2_20 (hash_out_2_20),
    .dout_valid_2_20 (hash_out_valid_2_20),
	.dout_2_21 (hash_out_2_21),
    .dout_valid_2_21 (hash_out_valid_2_21),
	.dout_2_22 (hash_out_2_22),
    .dout_valid_2_22 (hash_out_valid_2_22),
	.dout_2_23 (hash_out_2_23),
    .dout_valid_2_23 (hash_out_valid_2_23),
	.dout_2_24 (hash_out_2_24),
    .dout_valid_2_24 (hash_out_valid_2_24),
	.dout_2_25 (hash_out_2_25),
    .dout_valid_2_25 (hash_out_valid_2_25),
	.dout_2_26 (hash_out_2_26),
    .dout_valid_2_26 (hash_out_valid_2_26),
	.dout_2_27 (hash_out_2_27),
    .dout_valid_2_27 (hash_out_valid_2_27),
	.dout_2_28 (hash_out_2_28),
    .dout_valid_2_28 (hash_out_valid_2_28),
	.dout_2_29 (hash_out_2_29),
    .dout_valid_2_29 (hash_out_valid_2_29),
	.dout_2_30 (hash_out_2_30),
    .dout_valid_2_30 (hash_out_valid_2_30),
	.dout_2_31 (hash_out_2_31),
    .dout_valid_2_31 (hash_out_valid_2_31),
	.dout_3_0 (hash_out_3_0),
    .dout_valid_3_0 (hash_out_valid_3_0),
	.dout_3_1 (hash_out_3_1),
    .dout_valid_3_1 (hash_out_valid_3_1),
	.dout_3_2 (hash_out_3_2),
    .dout_valid_3_2 (hash_out_valid_3_2),
	.dout_3_3 (hash_out_3_3),
    .dout_valid_3_3 (hash_out_valid_3_3),
	.dout_3_4 (hash_out_3_4),
    .dout_valid_3_4 (hash_out_valid_3_4),
	.dout_3_5 (hash_out_3_5),
    .dout_valid_3_5 (hash_out_valid_3_5),
	.dout_3_6 (hash_out_3_6),
    .dout_valid_3_6 (hash_out_valid_3_6),
	.dout_3_7 (hash_out_3_7),
    .dout_valid_3_7 (hash_out_valid_3_7),
	.dout_3_8 (hash_out_3_8),
    .dout_valid_3_8 (hash_out_valid_3_8),
	.dout_3_9 (hash_out_3_9),
    .dout_valid_3_9 (hash_out_valid_3_9),
	.dout_3_10 (hash_out_3_10),
    .dout_valid_3_10 (hash_out_valid_3_10),
	.dout_3_11 (hash_out_3_11),
    .dout_valid_3_11 (hash_out_valid_3_11),
	.dout_3_12 (hash_out_3_12),
    .dout_valid_3_12 (hash_out_valid_3_12),
	.dout_3_13 (hash_out_3_13),
    .dout_valid_3_13 (hash_out_valid_3_13),
	.dout_3_14 (hash_out_3_14),
    .dout_valid_3_14 (hash_out_valid_3_14),
	.dout_3_15 (hash_out_3_15),
    .dout_valid_3_15 (hash_out_valid_3_15),
	.dout_3_16 (hash_out_3_16),
    .dout_valid_3_16 (hash_out_valid_3_16),
	.dout_3_17 (hash_out_3_17),
    .dout_valid_3_17 (hash_out_valid_3_17),
	.dout_3_18 (hash_out_3_18),
    .dout_valid_3_18 (hash_out_valid_3_18),
	.dout_3_19 (hash_out_3_19),
    .dout_valid_3_19 (hash_out_valid_3_19),
	.dout_3_20 (hash_out_3_20),
    .dout_valid_3_20 (hash_out_valid_3_20),
	.dout_3_21 (hash_out_3_21),
    .dout_valid_3_21 (hash_out_valid_3_21),
	.dout_3_22 (hash_out_3_22),
    .dout_valid_3_22 (hash_out_valid_3_22),
	.dout_3_23 (hash_out_3_23),
    .dout_valid_3_23 (hash_out_valid_3_23),
	.dout_3_24 (hash_out_3_24),
    .dout_valid_3_24 (hash_out_valid_3_24),
	.dout_3_25 (hash_out_3_25),
    .dout_valid_3_25 (hash_out_valid_3_25),
	.dout_3_26 (hash_out_3_26),
    .dout_valid_3_26 (hash_out_valid_3_26),
	.dout_3_27 (hash_out_3_27),
    .dout_valid_3_27 (hash_out_valid_3_27),
	.dout_3_28 (hash_out_3_28),
    .dout_valid_3_28 (hash_out_valid_3_28),
	.dout_3_29 (hash_out_3_29),
    .dout_valid_3_29 (hash_out_valid_3_29),
	.dout_3_30 (hash_out_3_30),
    .dout_valid_3_30 (hash_out_valid_3_30),
	.dout_3_31 (hash_out_3_31),
    .dout_valid_3_31 (hash_out_valid_3_31),
	.dout_4_0 (hash_out_4_0),
    .dout_valid_4_0 (hash_out_valid_4_0),
	.dout_4_1 (hash_out_4_1),
    .dout_valid_4_1 (hash_out_valid_4_1),
	.dout_4_2 (hash_out_4_2),
    .dout_valid_4_2 (hash_out_valid_4_2),
	.dout_4_3 (hash_out_4_3),
    .dout_valid_4_3 (hash_out_valid_4_3),
	.dout_4_4 (hash_out_4_4),
    .dout_valid_4_4 (hash_out_valid_4_4),
	.dout_4_5 (hash_out_4_5),
    .dout_valid_4_5 (hash_out_valid_4_5),
	.dout_4_6 (hash_out_4_6),
    .dout_valid_4_6 (hash_out_valid_4_6),
	.dout_4_7 (hash_out_4_7),
    .dout_valid_4_7 (hash_out_valid_4_7),
	.dout_4_8 (hash_out_4_8),
    .dout_valid_4_8 (hash_out_valid_4_8),
	.dout_4_9 (hash_out_4_9),
    .dout_valid_4_9 (hash_out_valid_4_9),
	.dout_4_10 (hash_out_4_10),
    .dout_valid_4_10 (hash_out_valid_4_10),
	.dout_4_11 (hash_out_4_11),
    .dout_valid_4_11 (hash_out_valid_4_11),
	.dout_4_12 (hash_out_4_12),
    .dout_valid_4_12 (hash_out_valid_4_12),
	.dout_4_13 (hash_out_4_13),
    .dout_valid_4_13 (hash_out_valid_4_13),
	.dout_4_14 (hash_out_4_14),
    .dout_valid_4_14 (hash_out_valid_4_14),
	.dout_4_15 (hash_out_4_15),
    .dout_valid_4_15 (hash_out_valid_4_15),
	.dout_4_16 (hash_out_4_16),
    .dout_valid_4_16 (hash_out_valid_4_16),
	.dout_4_17 (hash_out_4_17),
    .dout_valid_4_17 (hash_out_valid_4_17),
	.dout_4_18 (hash_out_4_18),
    .dout_valid_4_18 (hash_out_valid_4_18),
	.dout_4_19 (hash_out_4_19),
    .dout_valid_4_19 (hash_out_valid_4_19),
	.dout_4_20 (hash_out_4_20),
    .dout_valid_4_20 (hash_out_valid_4_20),
	.dout_4_21 (hash_out_4_21),
    .dout_valid_4_21 (hash_out_valid_4_21),
	.dout_4_22 (hash_out_4_22),
    .dout_valid_4_22 (hash_out_valid_4_22),
	.dout_4_23 (hash_out_4_23),
    .dout_valid_4_23 (hash_out_valid_4_23),
	.dout_4_24 (hash_out_4_24),
    .dout_valid_4_24 (hash_out_valid_4_24),
	.dout_4_25 (hash_out_4_25),
    .dout_valid_4_25 (hash_out_valid_4_25),
	.dout_4_26 (hash_out_4_26),
    .dout_valid_4_26 (hash_out_valid_4_26),
	.dout_4_27 (hash_out_4_27),
    .dout_valid_4_27 (hash_out_valid_4_27),
	.dout_4_28 (hash_out_4_28),
    .dout_valid_4_28 (hash_out_valid_4_28),
	.dout_4_29 (hash_out_4_29),
    .dout_valid_4_29 (hash_out_valid_4_29),
	.dout_4_30 (hash_out_4_30),
    .dout_valid_4_30 (hash_out_valid_4_30),
	.dout_4_31 (hash_out_4_31),
    .dout_valid_4_31 (hash_out_valid_4_31),
	.dout_5_0 (hash_out_5_0),
    .dout_valid_5_0 (hash_out_valid_5_0),
	.dout_5_1 (hash_out_5_1),
    .dout_valid_5_1 (hash_out_valid_5_1),
	.dout_5_2 (hash_out_5_2),
    .dout_valid_5_2 (hash_out_valid_5_2),
	.dout_5_3 (hash_out_5_3),
    .dout_valid_5_3 (hash_out_valid_5_3),
	.dout_5_4 (hash_out_5_4),
    .dout_valid_5_4 (hash_out_valid_5_4),
	.dout_5_5 (hash_out_5_5),
    .dout_valid_5_5 (hash_out_valid_5_5),
	.dout_5_6 (hash_out_5_6),
    .dout_valid_5_6 (hash_out_valid_5_6),
	.dout_5_7 (hash_out_5_7),
    .dout_valid_5_7 (hash_out_valid_5_7),
	.dout_5_8 (hash_out_5_8),
    .dout_valid_5_8 (hash_out_valid_5_8),
	.dout_5_9 (hash_out_5_9),
    .dout_valid_5_9 (hash_out_valid_5_9),
	.dout_5_10 (hash_out_5_10),
    .dout_valid_5_10 (hash_out_valid_5_10),
	.dout_5_11 (hash_out_5_11),
    .dout_valid_5_11 (hash_out_valid_5_11),
	.dout_5_12 (hash_out_5_12),
    .dout_valid_5_12 (hash_out_valid_5_12),
	.dout_5_13 (hash_out_5_13),
    .dout_valid_5_13 (hash_out_valid_5_13),
	.dout_5_14 (hash_out_5_14),
    .dout_valid_5_14 (hash_out_valid_5_14),
	.dout_5_15 (hash_out_5_15),
    .dout_valid_5_15 (hash_out_valid_5_15),
	.dout_5_16 (hash_out_5_16),
    .dout_valid_5_16 (hash_out_valid_5_16),
	.dout_5_17 (hash_out_5_17),
    .dout_valid_5_17 (hash_out_valid_5_17),
	.dout_5_18 (hash_out_5_18),
    .dout_valid_5_18 (hash_out_valid_5_18),
	.dout_5_19 (hash_out_5_19),
    .dout_valid_5_19 (hash_out_valid_5_19),
	.dout_5_20 (hash_out_5_20),
    .dout_valid_5_20 (hash_out_valid_5_20),
	.dout_5_21 (hash_out_5_21),
    .dout_valid_5_21 (hash_out_valid_5_21),
	.dout_5_22 (hash_out_5_22),
    .dout_valid_5_22 (hash_out_valid_5_22),
	.dout_5_23 (hash_out_5_23),
    .dout_valid_5_23 (hash_out_valid_5_23),
	.dout_5_24 (hash_out_5_24),
    .dout_valid_5_24 (hash_out_valid_5_24),
	.dout_5_25 (hash_out_5_25),
    .dout_valid_5_25 (hash_out_valid_5_25),
	.dout_5_26 (hash_out_5_26),
    .dout_valid_5_26 (hash_out_valid_5_26),
	.dout_5_27 (hash_out_5_27),
    .dout_valid_5_27 (hash_out_valid_5_27),
	.dout_5_28 (hash_out_5_28),
    .dout_valid_5_28 (hash_out_valid_5_28),
	.dout_5_29 (hash_out_5_29),
    .dout_valid_5_29 (hash_out_valid_5_29),
	.dout_5_30 (hash_out_5_30),
    .dout_valid_5_30 (hash_out_valid_5_30),
	.dout_5_31 (hash_out_5_31),
    .dout_valid_5_31 (hash_out_valid_5_31),
	.dout_6_0 (hash_out_6_0),
    .dout_valid_6_0 (hash_out_valid_6_0),
	.dout_6_1 (hash_out_6_1),
    .dout_valid_6_1 (hash_out_valid_6_1),
	.dout_6_2 (hash_out_6_2),
    .dout_valid_6_2 (hash_out_valid_6_2),
	.dout_6_3 (hash_out_6_3),
    .dout_valid_6_3 (hash_out_valid_6_3),
	.dout_6_4 (hash_out_6_4),
    .dout_valid_6_4 (hash_out_valid_6_4),
	.dout_6_5 (hash_out_6_5),
    .dout_valid_6_5 (hash_out_valid_6_5),
	.dout_6_6 (hash_out_6_6),
    .dout_valid_6_6 (hash_out_valid_6_6),
	.dout_6_7 (hash_out_6_7),
    .dout_valid_6_7 (hash_out_valid_6_7),
	.dout_6_8 (hash_out_6_8),
    .dout_valid_6_8 (hash_out_valid_6_8),
	.dout_6_9 (hash_out_6_9),
    .dout_valid_6_9 (hash_out_valid_6_9),
	.dout_6_10 (hash_out_6_10),
    .dout_valid_6_10 (hash_out_valid_6_10),
	.dout_6_11 (hash_out_6_11),
    .dout_valid_6_11 (hash_out_valid_6_11),
	.dout_6_12 (hash_out_6_12),
    .dout_valid_6_12 (hash_out_valid_6_12),
	.dout_6_13 (hash_out_6_13),
    .dout_valid_6_13 (hash_out_valid_6_13),
	.dout_6_14 (hash_out_6_14),
    .dout_valid_6_14 (hash_out_valid_6_14),
	.dout_6_15 (hash_out_6_15),
    .dout_valid_6_15 (hash_out_valid_6_15),
	.dout_6_16 (hash_out_6_16),
    .dout_valid_6_16 (hash_out_valid_6_16),
	.dout_6_17 (hash_out_6_17),
    .dout_valid_6_17 (hash_out_valid_6_17),
	.dout_6_18 (hash_out_6_18),
    .dout_valid_6_18 (hash_out_valid_6_18),
	.dout_6_19 (hash_out_6_19),
    .dout_valid_6_19 (hash_out_valid_6_19),
	.dout_6_20 (hash_out_6_20),
    .dout_valid_6_20 (hash_out_valid_6_20),
	.dout_6_21 (hash_out_6_21),
    .dout_valid_6_21 (hash_out_valid_6_21),
	.dout_6_22 (hash_out_6_22),
    .dout_valid_6_22 (hash_out_valid_6_22),
	.dout_6_23 (hash_out_6_23),
    .dout_valid_6_23 (hash_out_valid_6_23),
	.dout_6_24 (hash_out_6_24),
    .dout_valid_6_24 (hash_out_valid_6_24),
	.dout_6_25 (hash_out_6_25),
    .dout_valid_6_25 (hash_out_valid_6_25),
	.dout_6_26 (hash_out_6_26),
    .dout_valid_6_26 (hash_out_valid_6_26),
	.dout_6_27 (hash_out_6_27),
    .dout_valid_6_27 (hash_out_valid_6_27),
	.dout_6_28 (hash_out_6_28),
    .dout_valid_6_28 (hash_out_valid_6_28),
	.dout_6_29 (hash_out_6_29),
    .dout_valid_6_29 (hash_out_valid_6_29),
	.dout_6_30 (hash_out_6_30),
    .dout_valid_6_30 (hash_out_valid_6_30),
	.dout_6_31 (hash_out_6_31),
    .dout_valid_6_31 (hash_out_valid_6_31),
	.dout_7_0 (hash_out_7_0),
    .dout_valid_7_0 (hash_out_valid_7_0),
	.dout_7_1 (hash_out_7_1),
    .dout_valid_7_1 (hash_out_valid_7_1),
	.dout_7_2 (hash_out_7_2),
    .dout_valid_7_2 (hash_out_valid_7_2),
	.dout_7_3 (hash_out_7_3),
    .dout_valid_7_3 (hash_out_valid_7_3),
	.dout_7_4 (hash_out_7_4),
    .dout_valid_7_4 (hash_out_valid_7_4),
	.dout_7_5 (hash_out_7_5),
    .dout_valid_7_5 (hash_out_valid_7_5),
	.dout_7_6 (hash_out_7_6),
    .dout_valid_7_6 (hash_out_valid_7_6),
	.dout_7_7 (hash_out_7_7),
    .dout_valid_7_7 (hash_out_valid_7_7),
	.dout_7_8 (hash_out_7_8),
    .dout_valid_7_8 (hash_out_valid_7_8),
	.dout_7_9 (hash_out_7_9),
    .dout_valid_7_9 (hash_out_valid_7_9),
	.dout_7_10 (hash_out_7_10),
    .dout_valid_7_10 (hash_out_valid_7_10),
	.dout_7_11 (hash_out_7_11),
    .dout_valid_7_11 (hash_out_valid_7_11),
	.dout_7_12 (hash_out_7_12),
    .dout_valid_7_12 (hash_out_valid_7_12),
	.dout_7_13 (hash_out_7_13),
    .dout_valid_7_13 (hash_out_valid_7_13),
	.dout_7_14 (hash_out_7_14),
    .dout_valid_7_14 (hash_out_valid_7_14),
	.dout_7_15 (hash_out_7_15),
    .dout_valid_7_15 (hash_out_valid_7_15),
	.dout_7_16 (hash_out_7_16),
    .dout_valid_7_16 (hash_out_valid_7_16),
	.dout_7_17 (hash_out_7_17),
    .dout_valid_7_17 (hash_out_valid_7_17),
	.dout_7_18 (hash_out_7_18),
    .dout_valid_7_18 (hash_out_valid_7_18),
	.dout_7_19 (hash_out_7_19),
    .dout_valid_7_19 (hash_out_valid_7_19),
	.dout_7_20 (hash_out_7_20),
    .dout_valid_7_20 (hash_out_valid_7_20),
	.dout_7_21 (hash_out_7_21),
    .dout_valid_7_21 (hash_out_valid_7_21),
	.dout_7_22 (hash_out_7_22),
    .dout_valid_7_22 (hash_out_valid_7_22),
	.dout_7_23 (hash_out_7_23),
    .dout_valid_7_23 (hash_out_valid_7_23),
	.dout_7_24 (hash_out_7_24),
    .dout_valid_7_24 (hash_out_valid_7_24),
	.dout_7_25 (hash_out_7_25),
    .dout_valid_7_25 (hash_out_valid_7_25),
	.dout_7_26 (hash_out_7_26),
    .dout_valid_7_26 (hash_out_valid_7_26),
	.dout_7_27 (hash_out_7_27),
    .dout_valid_7_27 (hash_out_valid_7_27),
	.dout_7_28 (hash_out_7_28),
    .dout_valid_7_28 (hash_out_valid_7_28),
	.dout_7_29 (hash_out_7_29),
    .dout_valid_7_29 (hash_out_valid_7_29),
	.dout_7_30 (hash_out_7_30),
    .dout_valid_7_30 (hash_out_valid_7_30),
	.dout_7_31 (hash_out_7_31),
    .dout_valid_7_31 (hash_out_valid_7_31),
    .din (hash_in),
    .din_valid (hash_in_valid)
);

//Debug
/*
always@(*)begin
if(hash_out_valid_filter_0_0)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,0,hash_out_0_0);
end
if(hash_out_valid_filter_0_1)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,1,hash_out_0_1);
end
if(hash_out_valid_filter_0_2)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,2,hash_out_0_2);
end
if(hash_out_valid_filter_0_3)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,3,hash_out_0_3);
end
if(hash_out_valid_filter_0_4)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,4,hash_out_0_4);
end
if(hash_out_valid_filter_0_5)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,5,hash_out_0_5);
end
if(hash_out_valid_filter_0_6)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,6,hash_out_0_6);
end
if(hash_out_valid_filter_0_7)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,7,hash_out_0_7);
end
if(hash_out_valid_filter_0_8)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,8,hash_out_0_8);
end
if(hash_out_valid_filter_0_9)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,9,hash_out_0_9);
end
if(hash_out_valid_filter_0_10)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,10,hash_out_0_10);
end
if(hash_out_valid_filter_0_11)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,11,hash_out_0_11);
end
if(hash_out_valid_filter_0_12)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,12,hash_out_0_12);
end
if(hash_out_valid_filter_0_13)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,13,hash_out_0_13);
end
if(hash_out_valid_filter_0_14)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,14,hash_out_0_14);
end
if(hash_out_valid_filter_0_15)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,15,hash_out_0_15);
end
if(hash_out_valid_filter_0_16)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,16,hash_out_0_16);
end
if(hash_out_valid_filter_0_17)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,17,hash_out_0_17);
end
if(hash_out_valid_filter_0_18)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,18,hash_out_0_18);
end
if(hash_out_valid_filter_0_19)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,19,hash_out_0_19);
end
if(hash_out_valid_filter_0_20)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,20,hash_out_0_20);
end
if(hash_out_valid_filter_0_21)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,21,hash_out_0_21);
end
if(hash_out_valid_filter_0_22)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,22,hash_out_0_22);
end
if(hash_out_valid_filter_0_23)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,23,hash_out_0_23);
end
if(hash_out_valid_filter_0_24)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,24,hash_out_0_24);
end
if(hash_out_valid_filter_0_25)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,25,hash_out_0_25);
end
if(hash_out_valid_filter_0_26)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,26,hash_out_0_26);
end
if(hash_out_valid_filter_0_27)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,27,hash_out_0_27);
end
if(hash_out_valid_filter_0_28)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,28,hash_out_0_28);
end
if(hash_out_valid_filter_0_29)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,29,hash_out_0_29);
end
if(hash_out_valid_filter_0_30)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,30,hash_out_0_30);
end
if(hash_out_valid_filter_0_31)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        0,31,hash_out_0_31);
end
if(hash_out_valid_filter_1_0)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,0,hash_out_1_0);
end
if(hash_out_valid_filter_1_1)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,1,hash_out_1_1);
end
if(hash_out_valid_filter_1_2)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,2,hash_out_1_2);
end
if(hash_out_valid_filter_1_3)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,3,hash_out_1_3);
end
if(hash_out_valid_filter_1_4)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,4,hash_out_1_4);
end
if(hash_out_valid_filter_1_5)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,5,hash_out_1_5);
end
if(hash_out_valid_filter_1_6)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,6,hash_out_1_6);
end
if(hash_out_valid_filter_1_7)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,7,hash_out_1_7);
end
if(hash_out_valid_filter_1_8)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,8,hash_out_1_8);
end
if(hash_out_valid_filter_1_9)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,9,hash_out_1_9);
end
if(hash_out_valid_filter_1_10)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,10,hash_out_1_10);
end
if(hash_out_valid_filter_1_11)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,11,hash_out_1_11);
end
if(hash_out_valid_filter_1_12)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,12,hash_out_1_12);
end
if(hash_out_valid_filter_1_13)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,13,hash_out_1_13);
end
if(hash_out_valid_filter_1_14)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,14,hash_out_1_14);
end
if(hash_out_valid_filter_1_15)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,15,hash_out_1_15);
end
if(hash_out_valid_filter_1_16)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,16,hash_out_1_16);
end
if(hash_out_valid_filter_1_17)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,17,hash_out_1_17);
end
if(hash_out_valid_filter_1_18)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,18,hash_out_1_18);
end
if(hash_out_valid_filter_1_19)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,19,hash_out_1_19);
end
if(hash_out_valid_filter_1_20)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,20,hash_out_1_20);
end
if(hash_out_valid_filter_1_21)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,21,hash_out_1_21);
end
if(hash_out_valid_filter_1_22)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,22,hash_out_1_22);
end
if(hash_out_valid_filter_1_23)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,23,hash_out_1_23);
end
if(hash_out_valid_filter_1_24)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,24,hash_out_1_24);
end
if(hash_out_valid_filter_1_25)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,25,hash_out_1_25);
end
if(hash_out_valid_filter_1_26)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,26,hash_out_1_26);
end
if(hash_out_valid_filter_1_27)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,27,hash_out_1_27);
end
if(hash_out_valid_filter_1_28)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,28,hash_out_1_28);
end
if(hash_out_valid_filter_1_29)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,29,hash_out_1_29);
end
if(hash_out_valid_filter_1_30)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,30,hash_out_1_30);
end
if(hash_out_valid_filter_1_31)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        1,31,hash_out_1_31);
end
if(hash_out_valid_filter_2_0)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,0,hash_out_2_0);
end
if(hash_out_valid_filter_2_1)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,1,hash_out_2_1);
end
if(hash_out_valid_filter_2_2)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,2,hash_out_2_2);
end
if(hash_out_valid_filter_2_3)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,3,hash_out_2_3);
end
if(hash_out_valid_filter_2_4)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,4,hash_out_2_4);
end
if(hash_out_valid_filter_2_5)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,5,hash_out_2_5);
end
if(hash_out_valid_filter_2_6)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,6,hash_out_2_6);
end
if(hash_out_valid_filter_2_7)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,7,hash_out_2_7);
end
if(hash_out_valid_filter_2_8)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,8,hash_out_2_8);
end
if(hash_out_valid_filter_2_9)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,9,hash_out_2_9);
end
if(hash_out_valid_filter_2_10)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,10,hash_out_2_10);
end
if(hash_out_valid_filter_2_11)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,11,hash_out_2_11);
end
if(hash_out_valid_filter_2_12)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,12,hash_out_2_12);
end
if(hash_out_valid_filter_2_13)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,13,hash_out_2_13);
end
if(hash_out_valid_filter_2_14)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,14,hash_out_2_14);
end
if(hash_out_valid_filter_2_15)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,15,hash_out_2_15);
end
if(hash_out_valid_filter_2_16)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,16,hash_out_2_16);
end
if(hash_out_valid_filter_2_17)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,17,hash_out_2_17);
end
if(hash_out_valid_filter_2_18)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,18,hash_out_2_18);
end
if(hash_out_valid_filter_2_19)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,19,hash_out_2_19);
end
if(hash_out_valid_filter_2_20)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,20,hash_out_2_20);
end
if(hash_out_valid_filter_2_21)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,21,hash_out_2_21);
end
if(hash_out_valid_filter_2_22)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,22,hash_out_2_22);
end
if(hash_out_valid_filter_2_23)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,23,hash_out_2_23);
end
if(hash_out_valid_filter_2_24)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,24,hash_out_2_24);
end
if(hash_out_valid_filter_2_25)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,25,hash_out_2_25);
end
if(hash_out_valid_filter_2_26)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,26,hash_out_2_26);
end
if(hash_out_valid_filter_2_27)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,27,hash_out_2_27);
end
if(hash_out_valid_filter_2_28)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,28,hash_out_2_28);
end
if(hash_out_valid_filter_2_29)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,29,hash_out_2_29);
end
if(hash_out_valid_filter_2_30)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,30,hash_out_2_30);
end
if(hash_out_valid_filter_2_31)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        2,31,hash_out_2_31);
end
if(hash_out_valid_filter_3_0)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,0,hash_out_3_0);
end
if(hash_out_valid_filter_3_1)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,1,hash_out_3_1);
end
if(hash_out_valid_filter_3_2)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,2,hash_out_3_2);
end
if(hash_out_valid_filter_3_3)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,3,hash_out_3_3);
end
if(hash_out_valid_filter_3_4)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,4,hash_out_3_4);
end
if(hash_out_valid_filter_3_5)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,5,hash_out_3_5);
end
if(hash_out_valid_filter_3_6)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,6,hash_out_3_6);
end
if(hash_out_valid_filter_3_7)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,7,hash_out_3_7);
end
if(hash_out_valid_filter_3_8)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,8,hash_out_3_8);
end
if(hash_out_valid_filter_3_9)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,9,hash_out_3_9);
end
if(hash_out_valid_filter_3_10)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,10,hash_out_3_10);
end
if(hash_out_valid_filter_3_11)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,11,hash_out_3_11);
end
if(hash_out_valid_filter_3_12)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,12,hash_out_3_12);
end
if(hash_out_valid_filter_3_13)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,13,hash_out_3_13);
end
if(hash_out_valid_filter_3_14)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,14,hash_out_3_14);
end
if(hash_out_valid_filter_3_15)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,15,hash_out_3_15);
end
if(hash_out_valid_filter_3_16)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,16,hash_out_3_16);
end
if(hash_out_valid_filter_3_17)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,17,hash_out_3_17);
end
if(hash_out_valid_filter_3_18)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,18,hash_out_3_18);
end
if(hash_out_valid_filter_3_19)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,19,hash_out_3_19);
end
if(hash_out_valid_filter_3_20)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,20,hash_out_3_20);
end
if(hash_out_valid_filter_3_21)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,21,hash_out_3_21);
end
if(hash_out_valid_filter_3_22)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,22,hash_out_3_22);
end
if(hash_out_valid_filter_3_23)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,23,hash_out_3_23);
end
if(hash_out_valid_filter_3_24)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,24,hash_out_3_24);
end
if(hash_out_valid_filter_3_25)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,25,hash_out_3_25);
end
if(hash_out_valid_filter_3_26)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,26,hash_out_3_26);
end
if(hash_out_valid_filter_3_27)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,27,hash_out_3_27);
end
if(hash_out_valid_filter_3_28)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,28,hash_out_3_28);
end
if(hash_out_valid_filter_3_29)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,29,hash_out_3_29);
end
if(hash_out_valid_filter_3_30)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,30,hash_out_3_30);
end
if(hash_out_valid_filter_3_31)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        3,31,hash_out_3_31);
end
if(hash_out_valid_filter_4_0)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,0,hash_out_4_0);
end
if(hash_out_valid_filter_4_1)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,1,hash_out_4_1);
end
if(hash_out_valid_filter_4_2)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,2,hash_out_4_2);
end
if(hash_out_valid_filter_4_3)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,3,hash_out_4_3);
end
if(hash_out_valid_filter_4_4)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,4,hash_out_4_4);
end
if(hash_out_valid_filter_4_5)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,5,hash_out_4_5);
end
if(hash_out_valid_filter_4_6)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,6,hash_out_4_6);
end
if(hash_out_valid_filter_4_7)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,7,hash_out_4_7);
end
if(hash_out_valid_filter_4_8)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,8,hash_out_4_8);
end
if(hash_out_valid_filter_4_9)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,9,hash_out_4_9);
end
if(hash_out_valid_filter_4_10)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,10,hash_out_4_10);
end
if(hash_out_valid_filter_4_11)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,11,hash_out_4_11);
end
if(hash_out_valid_filter_4_12)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,12,hash_out_4_12);
end
if(hash_out_valid_filter_4_13)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,13,hash_out_4_13);
end
if(hash_out_valid_filter_4_14)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,14,hash_out_4_14);
end
if(hash_out_valid_filter_4_15)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,15,hash_out_4_15);
end
if(hash_out_valid_filter_4_16)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,16,hash_out_4_16);
end
if(hash_out_valid_filter_4_17)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,17,hash_out_4_17);
end
if(hash_out_valid_filter_4_18)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,18,hash_out_4_18);
end
if(hash_out_valid_filter_4_19)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,19,hash_out_4_19);
end
if(hash_out_valid_filter_4_20)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,20,hash_out_4_20);
end
if(hash_out_valid_filter_4_21)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,21,hash_out_4_21);
end
if(hash_out_valid_filter_4_22)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,22,hash_out_4_22);
end
if(hash_out_valid_filter_4_23)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,23,hash_out_4_23);
end
if(hash_out_valid_filter_4_24)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,24,hash_out_4_24);
end
if(hash_out_valid_filter_4_25)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,25,hash_out_4_25);
end
if(hash_out_valid_filter_4_26)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,26,hash_out_4_26);
end
if(hash_out_valid_filter_4_27)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,27,hash_out_4_27);
end
if(hash_out_valid_filter_4_28)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,28,hash_out_4_28);
end
if(hash_out_valid_filter_4_29)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,29,hash_out_4_29);
end
if(hash_out_valid_filter_4_30)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,30,hash_out_4_30);
end
if(hash_out_valid_filter_4_31)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        4,31,hash_out_4_31);
end
if(hash_out_valid_filter_5_0)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,0,hash_out_5_0);
end
if(hash_out_valid_filter_5_1)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,1,hash_out_5_1);
end
if(hash_out_valid_filter_5_2)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,2,hash_out_5_2);
end
if(hash_out_valid_filter_5_3)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,3,hash_out_5_3);
end
if(hash_out_valid_filter_5_4)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,4,hash_out_5_4);
end
if(hash_out_valid_filter_5_5)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,5,hash_out_5_5);
end
if(hash_out_valid_filter_5_6)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,6,hash_out_5_6);
end
if(hash_out_valid_filter_5_7)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,7,hash_out_5_7);
end
if(hash_out_valid_filter_5_8)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,8,hash_out_5_8);
end
if(hash_out_valid_filter_5_9)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,9,hash_out_5_9);
end
if(hash_out_valid_filter_5_10)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,10,hash_out_5_10);
end
if(hash_out_valid_filter_5_11)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,11,hash_out_5_11);
end
if(hash_out_valid_filter_5_12)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,12,hash_out_5_12);
end
if(hash_out_valid_filter_5_13)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,13,hash_out_5_13);
end
if(hash_out_valid_filter_5_14)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,14,hash_out_5_14);
end
if(hash_out_valid_filter_5_15)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,15,hash_out_5_15);
end
if(hash_out_valid_filter_5_16)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,16,hash_out_5_16);
end
if(hash_out_valid_filter_5_17)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,17,hash_out_5_17);
end
if(hash_out_valid_filter_5_18)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,18,hash_out_5_18);
end
if(hash_out_valid_filter_5_19)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,19,hash_out_5_19);
end
if(hash_out_valid_filter_5_20)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,20,hash_out_5_20);
end
if(hash_out_valid_filter_5_21)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,21,hash_out_5_21);
end
if(hash_out_valid_filter_5_22)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,22,hash_out_5_22);
end
if(hash_out_valid_filter_5_23)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,23,hash_out_5_23);
end
if(hash_out_valid_filter_5_24)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,24,hash_out_5_24);
end
if(hash_out_valid_filter_5_25)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,25,hash_out_5_25);
end
if(hash_out_valid_filter_5_26)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,26,hash_out_5_26);
end
if(hash_out_valid_filter_5_27)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,27,hash_out_5_27);
end
if(hash_out_valid_filter_5_28)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,28,hash_out_5_28);
end
if(hash_out_valid_filter_5_29)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,29,hash_out_5_29);
end
if(hash_out_valid_filter_5_30)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,30,hash_out_5_30);
end
if(hash_out_valid_filter_5_31)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        5,31,hash_out_5_31);
end
if(hash_out_valid_filter_6_0)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,0,hash_out_6_0);
end
if(hash_out_valid_filter_6_1)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,1,hash_out_6_1);
end
if(hash_out_valid_filter_6_2)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,2,hash_out_6_2);
end
if(hash_out_valid_filter_6_3)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,3,hash_out_6_3);
end
if(hash_out_valid_filter_6_4)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,4,hash_out_6_4);
end
if(hash_out_valid_filter_6_5)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,5,hash_out_6_5);
end
if(hash_out_valid_filter_6_6)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,6,hash_out_6_6);
end
if(hash_out_valid_filter_6_7)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,7,hash_out_6_7);
end
if(hash_out_valid_filter_6_8)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,8,hash_out_6_8);
end
if(hash_out_valid_filter_6_9)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,9,hash_out_6_9);
end
if(hash_out_valid_filter_6_10)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,10,hash_out_6_10);
end
if(hash_out_valid_filter_6_11)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,11,hash_out_6_11);
end
if(hash_out_valid_filter_6_12)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,12,hash_out_6_12);
end
if(hash_out_valid_filter_6_13)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,13,hash_out_6_13);
end
if(hash_out_valid_filter_6_14)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,14,hash_out_6_14);
end
if(hash_out_valid_filter_6_15)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,15,hash_out_6_15);
end
if(hash_out_valid_filter_6_16)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,16,hash_out_6_16);
end
if(hash_out_valid_filter_6_17)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,17,hash_out_6_17);
end
if(hash_out_valid_filter_6_18)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,18,hash_out_6_18);
end
if(hash_out_valid_filter_6_19)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,19,hash_out_6_19);
end
if(hash_out_valid_filter_6_20)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,20,hash_out_6_20);
end
if(hash_out_valid_filter_6_21)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,21,hash_out_6_21);
end
if(hash_out_valid_filter_6_22)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,22,hash_out_6_22);
end
if(hash_out_valid_filter_6_23)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,23,hash_out_6_23);
end
if(hash_out_valid_filter_6_24)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,24,hash_out_6_24);
end
if(hash_out_valid_filter_6_25)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,25,hash_out_6_25);
end
if(hash_out_valid_filter_6_26)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,26,hash_out_6_26);
end
if(hash_out_valid_filter_6_27)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,27,hash_out_6_27);
end
if(hash_out_valid_filter_6_28)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,28,hash_out_6_28);
end
if(hash_out_valid_filter_6_29)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,29,hash_out_6_29);
end
if(hash_out_valid_filter_6_30)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,30,hash_out_6_30);
end
if(hash_out_valid_filter_6_31)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        6,31,hash_out_6_31);
end
if(hash_out_valid_filter_7_0)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,0,hash_out_7_0);
end
if(hash_out_valid_filter_7_1)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,1,hash_out_7_1);
end
if(hash_out_valid_filter_7_2)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,2,hash_out_7_2);
end
if(hash_out_valid_filter_7_3)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,3,hash_out_7_3);
end
if(hash_out_valid_filter_7_4)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,4,hash_out_7_4);
end
if(hash_out_valid_filter_7_5)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,5,hash_out_7_5);
end
if(hash_out_valid_filter_7_6)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,6,hash_out_7_6);
end
if(hash_out_valid_filter_7_7)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,7,hash_out_7_7);
end
if(hash_out_valid_filter_7_8)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,8,hash_out_7_8);
end
if(hash_out_valid_filter_7_9)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,9,hash_out_7_9);
end
if(hash_out_valid_filter_7_10)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,10,hash_out_7_10);
end
if(hash_out_valid_filter_7_11)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,11,hash_out_7_11);
end
if(hash_out_valid_filter_7_12)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,12,hash_out_7_12);
end
if(hash_out_valid_filter_7_13)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,13,hash_out_7_13);
end
if(hash_out_valid_filter_7_14)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,14,hash_out_7_14);
end
if(hash_out_valid_filter_7_15)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,15,hash_out_7_15);
end
if(hash_out_valid_filter_7_16)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,16,hash_out_7_16);
end
if(hash_out_valid_filter_7_17)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,17,hash_out_7_17);
end
if(hash_out_valid_filter_7_18)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,18,hash_out_7_18);
end
if(hash_out_valid_filter_7_19)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,19,hash_out_7_19);
end
if(hash_out_valid_filter_7_20)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,20,hash_out_7_20);
end
if(hash_out_valid_filter_7_21)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,21,hash_out_7_21);
end
if(hash_out_valid_filter_7_22)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,22,hash_out_7_22);
end
if(hash_out_valid_filter_7_23)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,23,hash_out_7_23);
end
if(hash_out_valid_filter_7_24)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,24,hash_out_7_24);
end
if(hash_out_valid_filter_7_25)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,25,hash_out_7_25);
end
if(hash_out_valid_filter_7_26)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,26,hash_out_7_26);
end
if(hash_out_valid_filter_7_27)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,27,hash_out_7_27);
end
if(hash_out_valid_filter_7_28)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,28,hash_out_7_28);
end
if(hash_out_valid_filter_7_29)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,29,hash_out_7_29);
end
if(hash_out_valid_filter_7_30)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,30,hash_out_7_30);
end
if(hash_out_valid_filter_7_31)begin
    $display("Match: bucket %d, byte_position %d, RuleID %d",
        7,31,hash_out_7_31);
end
end
*/
`endif
endmodule //top
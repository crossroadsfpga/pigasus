`include "./src/struct_s.sv"
//`define DUMMY
//`define DEBUG
module string_matcher (
    input  logic                 front_clk,
    input  logic                 front_rst,
    input  logic                 back_clk,
    input  logic                 back_rst,
    input  logic [FP_DWIDTH-1:0] in_pkt_data,
    input  logic                 in_pkt_valid,
    input  logic                 in_pkt_sop,
    input  logic                 in_pkt_eop,
    input  logic [FP_EWIDTH-1:0] in_pkt_empty,
    output logic                 in_pkt_ready,
    output logic [511:0]         out_usr_data,
    output logic                 out_usr_valid,
    output logic                 out_usr_sop,
    output logic                 out_usr_eop,
    output logic [5:0]           out_usr_empty,
    input  logic                 out_usr_ready
);

`ifdef DUMMY

assign in_pkt_ready = 1;
assign out_usr_data = 0;
assign out_usr_sop  = out_usr_eop;
assign out_usr_empty = 0;
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dummy_FIFO"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (0),
    .FULL_LEVEL       (20),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (META_WIDTH),
    .FIFO_DEPTH       (32)
) in_meta_fifo (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (1'b1),
    .in_valid          (in_pkt_valid & in_pkt_eop),
    .in_ready          (),
    .out_data          (out_usr_eop),
    .out_valid         (out_usr_valid),
    .out_ready         (out_usr_ready),
    .fill_level        (),
    .almost_full       (),
    .overflow          ()
);

`else
///////NOT DUMMY////////////
logic [FP_DWIDTH-1:0]  piped_pkt_data;
logic                  piped_pkt_valid;
logic                  piped_pkt_sop;
logic                  piped_pkt_eop;
logic [FP_EWIDTH-1:0]  piped_pkt_empty;
logic [FP_DWIDTH-1:0]  piped_pkt_data_swap;
logic                  piped_pkt_almost_full;

//debug
logic [31:0] in_pkt_cnt;
logic [31:0] out_rule_cnt;
logic [31:0] out_rule_last_cnt;


logic [RID_WIDTH-1:0] hash_out_0_0;
logic hash_out_valid_filter_0_0;
rule_s_t din_0_0;
rule_s_t din_0_0_r1;
rule_s_t din_0_0_r2;
logic din_valid_0_0;
logic din_valid_0_0_r1;
logic din_valid_0_0_r2;
logic din_ready_0_0;
logic din_almost_full_0_0;
logic [31:0] din_csr_readdata_0_0;
rule_s_t back_data_0_0;
logic    back_valid_0_0;
logic    back_ready_0_0;
logic [RID_WIDTH-1:0] hash_out_0_1;
logic hash_out_valid_filter_0_1;
rule_s_t din_0_1;
rule_s_t din_0_1_r1;
rule_s_t din_0_1_r2;
logic din_valid_0_1;
logic din_valid_0_1_r1;
logic din_valid_0_1_r2;
logic din_ready_0_1;
logic din_almost_full_0_1;
logic [31:0] din_csr_readdata_0_1;
rule_s_t back_data_0_1;
logic    back_valid_0_1;
logic    back_ready_0_1;
logic [RID_WIDTH-1:0] hash_out_0_2;
logic hash_out_valid_filter_0_2;
rule_s_t din_0_2;
rule_s_t din_0_2_r1;
rule_s_t din_0_2_r2;
logic din_valid_0_2;
logic din_valid_0_2_r1;
logic din_valid_0_2_r2;
logic din_ready_0_2;
logic din_almost_full_0_2;
logic [31:0] din_csr_readdata_0_2;
rule_s_t back_data_0_2;
logic    back_valid_0_2;
logic    back_ready_0_2;
logic [RID_WIDTH-1:0] hash_out_0_3;
logic hash_out_valid_filter_0_3;
rule_s_t din_0_3;
rule_s_t din_0_3_r1;
rule_s_t din_0_3_r2;
logic din_valid_0_3;
logic din_valid_0_3_r1;
logic din_valid_0_3_r2;
logic din_ready_0_3;
logic din_almost_full_0_3;
logic [31:0] din_csr_readdata_0_3;
rule_s_t back_data_0_3;
logic    back_valid_0_3;
logic    back_ready_0_3;
logic [RID_WIDTH-1:0] hash_out_0_4;
logic hash_out_valid_filter_0_4;
rule_s_t din_0_4;
rule_s_t din_0_4_r1;
rule_s_t din_0_4_r2;
logic din_valid_0_4;
logic din_valid_0_4_r1;
logic din_valid_0_4_r2;
logic din_ready_0_4;
logic din_almost_full_0_4;
logic [31:0] din_csr_readdata_0_4;
rule_s_t back_data_0_4;
logic    back_valid_0_4;
logic    back_ready_0_4;
logic [RID_WIDTH-1:0] hash_out_0_5;
logic hash_out_valid_filter_0_5;
rule_s_t din_0_5;
rule_s_t din_0_5_r1;
rule_s_t din_0_5_r2;
logic din_valid_0_5;
logic din_valid_0_5_r1;
logic din_valid_0_5_r2;
logic din_ready_0_5;
logic din_almost_full_0_5;
logic [31:0] din_csr_readdata_0_5;
rule_s_t back_data_0_5;
logic    back_valid_0_5;
logic    back_ready_0_5;
logic [RID_WIDTH-1:0] hash_out_0_6;
logic hash_out_valid_filter_0_6;
rule_s_t din_0_6;
rule_s_t din_0_6_r1;
rule_s_t din_0_6_r2;
logic din_valid_0_6;
logic din_valid_0_6_r1;
logic din_valid_0_6_r2;
logic din_ready_0_6;
logic din_almost_full_0_6;
logic [31:0] din_csr_readdata_0_6;
rule_s_t back_data_0_6;
logic    back_valid_0_6;
logic    back_ready_0_6;
logic [RID_WIDTH-1:0] hash_out_0_7;
logic hash_out_valid_filter_0_7;
rule_s_t din_0_7;
rule_s_t din_0_7_r1;
rule_s_t din_0_7_r2;
logic din_valid_0_7;
logic din_valid_0_7_r1;
logic din_valid_0_7_r2;
logic din_ready_0_7;
logic din_almost_full_0_7;
logic [31:0] din_csr_readdata_0_7;
rule_s_t back_data_0_7;
logic    back_valid_0_7;
logic    back_ready_0_7;
logic [RID_WIDTH-1:0] hash_out_0_8;
logic hash_out_valid_filter_0_8;
rule_s_t din_0_8;
rule_s_t din_0_8_r1;
rule_s_t din_0_8_r2;
logic din_valid_0_8;
logic din_valid_0_8_r1;
logic din_valid_0_8_r2;
logic din_ready_0_8;
logic din_almost_full_0_8;
logic [31:0] din_csr_readdata_0_8;
rule_s_t back_data_0_8;
logic    back_valid_0_8;
logic    back_ready_0_8;
logic [RID_WIDTH-1:0] hash_out_0_9;
logic hash_out_valid_filter_0_9;
rule_s_t din_0_9;
rule_s_t din_0_9_r1;
rule_s_t din_0_9_r2;
logic din_valid_0_9;
logic din_valid_0_9_r1;
logic din_valid_0_9_r2;
logic din_ready_0_9;
logic din_almost_full_0_9;
logic [31:0] din_csr_readdata_0_9;
rule_s_t back_data_0_9;
logic    back_valid_0_9;
logic    back_ready_0_9;
logic [RID_WIDTH-1:0] hash_out_0_10;
logic hash_out_valid_filter_0_10;
rule_s_t din_0_10;
rule_s_t din_0_10_r1;
rule_s_t din_0_10_r2;
logic din_valid_0_10;
logic din_valid_0_10_r1;
logic din_valid_0_10_r2;
logic din_ready_0_10;
logic din_almost_full_0_10;
logic [31:0] din_csr_readdata_0_10;
rule_s_t back_data_0_10;
logic    back_valid_0_10;
logic    back_ready_0_10;
logic [RID_WIDTH-1:0] hash_out_0_11;
logic hash_out_valid_filter_0_11;
rule_s_t din_0_11;
rule_s_t din_0_11_r1;
rule_s_t din_0_11_r2;
logic din_valid_0_11;
logic din_valid_0_11_r1;
logic din_valid_0_11_r2;
logic din_ready_0_11;
logic din_almost_full_0_11;
logic [31:0] din_csr_readdata_0_11;
rule_s_t back_data_0_11;
logic    back_valid_0_11;
logic    back_ready_0_11;
logic [RID_WIDTH-1:0] hash_out_0_12;
logic hash_out_valid_filter_0_12;
rule_s_t din_0_12;
rule_s_t din_0_12_r1;
rule_s_t din_0_12_r2;
logic din_valid_0_12;
logic din_valid_0_12_r1;
logic din_valid_0_12_r2;
logic din_ready_0_12;
logic din_almost_full_0_12;
logic [31:0] din_csr_readdata_0_12;
rule_s_t back_data_0_12;
logic    back_valid_0_12;
logic    back_ready_0_12;
logic [RID_WIDTH-1:0] hash_out_0_13;
logic hash_out_valid_filter_0_13;
rule_s_t din_0_13;
rule_s_t din_0_13_r1;
rule_s_t din_0_13_r2;
logic din_valid_0_13;
logic din_valid_0_13_r1;
logic din_valid_0_13_r2;
logic din_ready_0_13;
logic din_almost_full_0_13;
logic [31:0] din_csr_readdata_0_13;
rule_s_t back_data_0_13;
logic    back_valid_0_13;
logic    back_ready_0_13;
logic [RID_WIDTH-1:0] hash_out_0_14;
logic hash_out_valid_filter_0_14;
rule_s_t din_0_14;
rule_s_t din_0_14_r1;
rule_s_t din_0_14_r2;
logic din_valid_0_14;
logic din_valid_0_14_r1;
logic din_valid_0_14_r2;
logic din_ready_0_14;
logic din_almost_full_0_14;
logic [31:0] din_csr_readdata_0_14;
rule_s_t back_data_0_14;
logic    back_valid_0_14;
logic    back_ready_0_14;
logic [RID_WIDTH-1:0] hash_out_0_15;
logic hash_out_valid_filter_0_15;
rule_s_t din_0_15;
rule_s_t din_0_15_r1;
rule_s_t din_0_15_r2;
logic din_valid_0_15;
logic din_valid_0_15_r1;
logic din_valid_0_15_r2;
logic din_ready_0_15;
logic din_almost_full_0_15;
logic [31:0] din_csr_readdata_0_15;
rule_s_t back_data_0_15;
logic    back_valid_0_15;
logic    back_ready_0_15;
logic [RID_WIDTH-1:0] hash_out_0_16;
logic hash_out_valid_filter_0_16;
rule_s_t din_0_16;
rule_s_t din_0_16_r1;
rule_s_t din_0_16_r2;
logic din_valid_0_16;
logic din_valid_0_16_r1;
logic din_valid_0_16_r2;
logic din_ready_0_16;
logic din_almost_full_0_16;
logic [31:0] din_csr_readdata_0_16;
rule_s_t back_data_0_16;
logic    back_valid_0_16;
logic    back_ready_0_16;
logic [RID_WIDTH-1:0] hash_out_0_17;
logic hash_out_valid_filter_0_17;
rule_s_t din_0_17;
rule_s_t din_0_17_r1;
rule_s_t din_0_17_r2;
logic din_valid_0_17;
logic din_valid_0_17_r1;
logic din_valid_0_17_r2;
logic din_ready_0_17;
logic din_almost_full_0_17;
logic [31:0] din_csr_readdata_0_17;
rule_s_t back_data_0_17;
logic    back_valid_0_17;
logic    back_ready_0_17;
logic [RID_WIDTH-1:0] hash_out_0_18;
logic hash_out_valid_filter_0_18;
rule_s_t din_0_18;
rule_s_t din_0_18_r1;
rule_s_t din_0_18_r2;
logic din_valid_0_18;
logic din_valid_0_18_r1;
logic din_valid_0_18_r2;
logic din_ready_0_18;
logic din_almost_full_0_18;
logic [31:0] din_csr_readdata_0_18;
rule_s_t back_data_0_18;
logic    back_valid_0_18;
logic    back_ready_0_18;
logic [RID_WIDTH-1:0] hash_out_0_19;
logic hash_out_valid_filter_0_19;
rule_s_t din_0_19;
rule_s_t din_0_19_r1;
rule_s_t din_0_19_r2;
logic din_valid_0_19;
logic din_valid_0_19_r1;
logic din_valid_0_19_r2;
logic din_ready_0_19;
logic din_almost_full_0_19;
logic [31:0] din_csr_readdata_0_19;
rule_s_t back_data_0_19;
logic    back_valid_0_19;
logic    back_ready_0_19;
logic [RID_WIDTH-1:0] hash_out_0_20;
logic hash_out_valid_filter_0_20;
rule_s_t din_0_20;
rule_s_t din_0_20_r1;
rule_s_t din_0_20_r2;
logic din_valid_0_20;
logic din_valid_0_20_r1;
logic din_valid_0_20_r2;
logic din_ready_0_20;
logic din_almost_full_0_20;
logic [31:0] din_csr_readdata_0_20;
rule_s_t back_data_0_20;
logic    back_valid_0_20;
logic    back_ready_0_20;
logic [RID_WIDTH-1:0] hash_out_0_21;
logic hash_out_valid_filter_0_21;
rule_s_t din_0_21;
rule_s_t din_0_21_r1;
rule_s_t din_0_21_r2;
logic din_valid_0_21;
logic din_valid_0_21_r1;
logic din_valid_0_21_r2;
logic din_ready_0_21;
logic din_almost_full_0_21;
logic [31:0] din_csr_readdata_0_21;
rule_s_t back_data_0_21;
logic    back_valid_0_21;
logic    back_ready_0_21;
logic [RID_WIDTH-1:0] hash_out_0_22;
logic hash_out_valid_filter_0_22;
rule_s_t din_0_22;
rule_s_t din_0_22_r1;
rule_s_t din_0_22_r2;
logic din_valid_0_22;
logic din_valid_0_22_r1;
logic din_valid_0_22_r2;
logic din_ready_0_22;
logic din_almost_full_0_22;
logic [31:0] din_csr_readdata_0_22;
rule_s_t back_data_0_22;
logic    back_valid_0_22;
logic    back_ready_0_22;
logic [RID_WIDTH-1:0] hash_out_0_23;
logic hash_out_valid_filter_0_23;
rule_s_t din_0_23;
rule_s_t din_0_23_r1;
rule_s_t din_0_23_r2;
logic din_valid_0_23;
logic din_valid_0_23_r1;
logic din_valid_0_23_r2;
logic din_ready_0_23;
logic din_almost_full_0_23;
logic [31:0] din_csr_readdata_0_23;
rule_s_t back_data_0_23;
logic    back_valid_0_23;
logic    back_ready_0_23;
logic [RID_WIDTH-1:0] hash_out_0_24;
logic hash_out_valid_filter_0_24;
rule_s_t din_0_24;
rule_s_t din_0_24_r1;
rule_s_t din_0_24_r2;
logic din_valid_0_24;
logic din_valid_0_24_r1;
logic din_valid_0_24_r2;
logic din_ready_0_24;
logic din_almost_full_0_24;
logic [31:0] din_csr_readdata_0_24;
rule_s_t back_data_0_24;
logic    back_valid_0_24;
logic    back_ready_0_24;
logic [RID_WIDTH-1:0] hash_out_0_25;
logic hash_out_valid_filter_0_25;
rule_s_t din_0_25;
rule_s_t din_0_25_r1;
rule_s_t din_0_25_r2;
logic din_valid_0_25;
logic din_valid_0_25_r1;
logic din_valid_0_25_r2;
logic din_ready_0_25;
logic din_almost_full_0_25;
logic [31:0] din_csr_readdata_0_25;
rule_s_t back_data_0_25;
logic    back_valid_0_25;
logic    back_ready_0_25;
logic [RID_WIDTH-1:0] hash_out_0_26;
logic hash_out_valid_filter_0_26;
rule_s_t din_0_26;
rule_s_t din_0_26_r1;
rule_s_t din_0_26_r2;
logic din_valid_0_26;
logic din_valid_0_26_r1;
logic din_valid_0_26_r2;
logic din_ready_0_26;
logic din_almost_full_0_26;
logic [31:0] din_csr_readdata_0_26;
rule_s_t back_data_0_26;
logic    back_valid_0_26;
logic    back_ready_0_26;
logic [RID_WIDTH-1:0] hash_out_0_27;
logic hash_out_valid_filter_0_27;
rule_s_t din_0_27;
rule_s_t din_0_27_r1;
rule_s_t din_0_27_r2;
logic din_valid_0_27;
logic din_valid_0_27_r1;
logic din_valid_0_27_r2;
logic din_ready_0_27;
logic din_almost_full_0_27;
logic [31:0] din_csr_readdata_0_27;
rule_s_t back_data_0_27;
logic    back_valid_0_27;
logic    back_ready_0_27;
logic [RID_WIDTH-1:0] hash_out_0_28;
logic hash_out_valid_filter_0_28;
rule_s_t din_0_28;
rule_s_t din_0_28_r1;
rule_s_t din_0_28_r2;
logic din_valid_0_28;
logic din_valid_0_28_r1;
logic din_valid_0_28_r2;
logic din_ready_0_28;
logic din_almost_full_0_28;
logic [31:0] din_csr_readdata_0_28;
rule_s_t back_data_0_28;
logic    back_valid_0_28;
logic    back_ready_0_28;
logic [RID_WIDTH-1:0] hash_out_0_29;
logic hash_out_valid_filter_0_29;
rule_s_t din_0_29;
rule_s_t din_0_29_r1;
rule_s_t din_0_29_r2;
logic din_valid_0_29;
logic din_valid_0_29_r1;
logic din_valid_0_29_r2;
logic din_ready_0_29;
logic din_almost_full_0_29;
logic [31:0] din_csr_readdata_0_29;
rule_s_t back_data_0_29;
logic    back_valid_0_29;
logic    back_ready_0_29;
logic [RID_WIDTH-1:0] hash_out_0_30;
logic hash_out_valid_filter_0_30;
rule_s_t din_0_30;
rule_s_t din_0_30_r1;
rule_s_t din_0_30_r2;
logic din_valid_0_30;
logic din_valid_0_30_r1;
logic din_valid_0_30_r2;
logic din_ready_0_30;
logic din_almost_full_0_30;
logic [31:0] din_csr_readdata_0_30;
rule_s_t back_data_0_30;
logic    back_valid_0_30;
logic    back_ready_0_30;
logic [RID_WIDTH-1:0] hash_out_0_31;
logic hash_out_valid_filter_0_31;
rule_s_t din_0_31;
rule_s_t din_0_31_r1;
rule_s_t din_0_31_r2;
logic din_valid_0_31;
logic din_valid_0_31_r1;
logic din_valid_0_31_r2;
logic din_ready_0_31;
logic din_almost_full_0_31;
logic [31:0] din_csr_readdata_0_31;
rule_s_t back_data_0_31;
logic    back_valid_0_31;
logic    back_ready_0_31;
logic [RID_WIDTH-1:0] hash_out_1_0;
logic hash_out_valid_filter_1_0;
rule_s_t din_1_0;
rule_s_t din_1_0_r1;
rule_s_t din_1_0_r2;
logic din_valid_1_0;
logic din_valid_1_0_r1;
logic din_valid_1_0_r2;
logic din_ready_1_0;
logic din_almost_full_1_0;
logic [31:0] din_csr_readdata_1_0;
rule_s_t back_data_1_0;
logic    back_valid_1_0;
logic    back_ready_1_0;
logic [RID_WIDTH-1:0] hash_out_1_1;
logic hash_out_valid_filter_1_1;
rule_s_t din_1_1;
rule_s_t din_1_1_r1;
rule_s_t din_1_1_r2;
logic din_valid_1_1;
logic din_valid_1_1_r1;
logic din_valid_1_1_r2;
logic din_ready_1_1;
logic din_almost_full_1_1;
logic [31:0] din_csr_readdata_1_1;
rule_s_t back_data_1_1;
logic    back_valid_1_1;
logic    back_ready_1_1;
logic [RID_WIDTH-1:0] hash_out_1_2;
logic hash_out_valid_filter_1_2;
rule_s_t din_1_2;
rule_s_t din_1_2_r1;
rule_s_t din_1_2_r2;
logic din_valid_1_2;
logic din_valid_1_2_r1;
logic din_valid_1_2_r2;
logic din_ready_1_2;
logic din_almost_full_1_2;
logic [31:0] din_csr_readdata_1_2;
rule_s_t back_data_1_2;
logic    back_valid_1_2;
logic    back_ready_1_2;
logic [RID_WIDTH-1:0] hash_out_1_3;
logic hash_out_valid_filter_1_3;
rule_s_t din_1_3;
rule_s_t din_1_3_r1;
rule_s_t din_1_3_r2;
logic din_valid_1_3;
logic din_valid_1_3_r1;
logic din_valid_1_3_r2;
logic din_ready_1_3;
logic din_almost_full_1_3;
logic [31:0] din_csr_readdata_1_3;
rule_s_t back_data_1_3;
logic    back_valid_1_3;
logic    back_ready_1_3;
logic [RID_WIDTH-1:0] hash_out_1_4;
logic hash_out_valid_filter_1_4;
rule_s_t din_1_4;
rule_s_t din_1_4_r1;
rule_s_t din_1_4_r2;
logic din_valid_1_4;
logic din_valid_1_4_r1;
logic din_valid_1_4_r2;
logic din_ready_1_4;
logic din_almost_full_1_4;
logic [31:0] din_csr_readdata_1_4;
rule_s_t back_data_1_4;
logic    back_valid_1_4;
logic    back_ready_1_4;
logic [RID_WIDTH-1:0] hash_out_1_5;
logic hash_out_valid_filter_1_5;
rule_s_t din_1_5;
rule_s_t din_1_5_r1;
rule_s_t din_1_5_r2;
logic din_valid_1_5;
logic din_valid_1_5_r1;
logic din_valid_1_5_r2;
logic din_ready_1_5;
logic din_almost_full_1_5;
logic [31:0] din_csr_readdata_1_5;
rule_s_t back_data_1_5;
logic    back_valid_1_5;
logic    back_ready_1_5;
logic [RID_WIDTH-1:0] hash_out_1_6;
logic hash_out_valid_filter_1_6;
rule_s_t din_1_6;
rule_s_t din_1_6_r1;
rule_s_t din_1_6_r2;
logic din_valid_1_6;
logic din_valid_1_6_r1;
logic din_valid_1_6_r2;
logic din_ready_1_6;
logic din_almost_full_1_6;
logic [31:0] din_csr_readdata_1_6;
rule_s_t back_data_1_6;
logic    back_valid_1_6;
logic    back_ready_1_6;
logic [RID_WIDTH-1:0] hash_out_1_7;
logic hash_out_valid_filter_1_7;
rule_s_t din_1_7;
rule_s_t din_1_7_r1;
rule_s_t din_1_7_r2;
logic din_valid_1_7;
logic din_valid_1_7_r1;
logic din_valid_1_7_r2;
logic din_ready_1_7;
logic din_almost_full_1_7;
logic [31:0] din_csr_readdata_1_7;
rule_s_t back_data_1_7;
logic    back_valid_1_7;
logic    back_ready_1_7;
logic [RID_WIDTH-1:0] hash_out_1_8;
logic hash_out_valid_filter_1_8;
rule_s_t din_1_8;
rule_s_t din_1_8_r1;
rule_s_t din_1_8_r2;
logic din_valid_1_8;
logic din_valid_1_8_r1;
logic din_valid_1_8_r2;
logic din_ready_1_8;
logic din_almost_full_1_8;
logic [31:0] din_csr_readdata_1_8;
rule_s_t back_data_1_8;
logic    back_valid_1_8;
logic    back_ready_1_8;
logic [RID_WIDTH-1:0] hash_out_1_9;
logic hash_out_valid_filter_1_9;
rule_s_t din_1_9;
rule_s_t din_1_9_r1;
rule_s_t din_1_9_r2;
logic din_valid_1_9;
logic din_valid_1_9_r1;
logic din_valid_1_9_r2;
logic din_ready_1_9;
logic din_almost_full_1_9;
logic [31:0] din_csr_readdata_1_9;
rule_s_t back_data_1_9;
logic    back_valid_1_9;
logic    back_ready_1_9;
logic [RID_WIDTH-1:0] hash_out_1_10;
logic hash_out_valid_filter_1_10;
rule_s_t din_1_10;
rule_s_t din_1_10_r1;
rule_s_t din_1_10_r2;
logic din_valid_1_10;
logic din_valid_1_10_r1;
logic din_valid_1_10_r2;
logic din_ready_1_10;
logic din_almost_full_1_10;
logic [31:0] din_csr_readdata_1_10;
rule_s_t back_data_1_10;
logic    back_valid_1_10;
logic    back_ready_1_10;
logic [RID_WIDTH-1:0] hash_out_1_11;
logic hash_out_valid_filter_1_11;
rule_s_t din_1_11;
rule_s_t din_1_11_r1;
rule_s_t din_1_11_r2;
logic din_valid_1_11;
logic din_valid_1_11_r1;
logic din_valid_1_11_r2;
logic din_ready_1_11;
logic din_almost_full_1_11;
logic [31:0] din_csr_readdata_1_11;
rule_s_t back_data_1_11;
logic    back_valid_1_11;
logic    back_ready_1_11;
logic [RID_WIDTH-1:0] hash_out_1_12;
logic hash_out_valid_filter_1_12;
rule_s_t din_1_12;
rule_s_t din_1_12_r1;
rule_s_t din_1_12_r2;
logic din_valid_1_12;
logic din_valid_1_12_r1;
logic din_valid_1_12_r2;
logic din_ready_1_12;
logic din_almost_full_1_12;
logic [31:0] din_csr_readdata_1_12;
rule_s_t back_data_1_12;
logic    back_valid_1_12;
logic    back_ready_1_12;
logic [RID_WIDTH-1:0] hash_out_1_13;
logic hash_out_valid_filter_1_13;
rule_s_t din_1_13;
rule_s_t din_1_13_r1;
rule_s_t din_1_13_r2;
logic din_valid_1_13;
logic din_valid_1_13_r1;
logic din_valid_1_13_r2;
logic din_ready_1_13;
logic din_almost_full_1_13;
logic [31:0] din_csr_readdata_1_13;
rule_s_t back_data_1_13;
logic    back_valid_1_13;
logic    back_ready_1_13;
logic [RID_WIDTH-1:0] hash_out_1_14;
logic hash_out_valid_filter_1_14;
rule_s_t din_1_14;
rule_s_t din_1_14_r1;
rule_s_t din_1_14_r2;
logic din_valid_1_14;
logic din_valid_1_14_r1;
logic din_valid_1_14_r2;
logic din_ready_1_14;
logic din_almost_full_1_14;
logic [31:0] din_csr_readdata_1_14;
rule_s_t back_data_1_14;
logic    back_valid_1_14;
logic    back_ready_1_14;
logic [RID_WIDTH-1:0] hash_out_1_15;
logic hash_out_valid_filter_1_15;
rule_s_t din_1_15;
rule_s_t din_1_15_r1;
rule_s_t din_1_15_r2;
logic din_valid_1_15;
logic din_valid_1_15_r1;
logic din_valid_1_15_r2;
logic din_ready_1_15;
logic din_almost_full_1_15;
logic [31:0] din_csr_readdata_1_15;
rule_s_t back_data_1_15;
logic    back_valid_1_15;
logic    back_ready_1_15;
logic [RID_WIDTH-1:0] hash_out_1_16;
logic hash_out_valid_filter_1_16;
rule_s_t din_1_16;
rule_s_t din_1_16_r1;
rule_s_t din_1_16_r2;
logic din_valid_1_16;
logic din_valid_1_16_r1;
logic din_valid_1_16_r2;
logic din_ready_1_16;
logic din_almost_full_1_16;
logic [31:0] din_csr_readdata_1_16;
rule_s_t back_data_1_16;
logic    back_valid_1_16;
logic    back_ready_1_16;
logic [RID_WIDTH-1:0] hash_out_1_17;
logic hash_out_valid_filter_1_17;
rule_s_t din_1_17;
rule_s_t din_1_17_r1;
rule_s_t din_1_17_r2;
logic din_valid_1_17;
logic din_valid_1_17_r1;
logic din_valid_1_17_r2;
logic din_ready_1_17;
logic din_almost_full_1_17;
logic [31:0] din_csr_readdata_1_17;
rule_s_t back_data_1_17;
logic    back_valid_1_17;
logic    back_ready_1_17;
logic [RID_WIDTH-1:0] hash_out_1_18;
logic hash_out_valid_filter_1_18;
rule_s_t din_1_18;
rule_s_t din_1_18_r1;
rule_s_t din_1_18_r2;
logic din_valid_1_18;
logic din_valid_1_18_r1;
logic din_valid_1_18_r2;
logic din_ready_1_18;
logic din_almost_full_1_18;
logic [31:0] din_csr_readdata_1_18;
rule_s_t back_data_1_18;
logic    back_valid_1_18;
logic    back_ready_1_18;
logic [RID_WIDTH-1:0] hash_out_1_19;
logic hash_out_valid_filter_1_19;
rule_s_t din_1_19;
rule_s_t din_1_19_r1;
rule_s_t din_1_19_r2;
logic din_valid_1_19;
logic din_valid_1_19_r1;
logic din_valid_1_19_r2;
logic din_ready_1_19;
logic din_almost_full_1_19;
logic [31:0] din_csr_readdata_1_19;
rule_s_t back_data_1_19;
logic    back_valid_1_19;
logic    back_ready_1_19;
logic [RID_WIDTH-1:0] hash_out_1_20;
logic hash_out_valid_filter_1_20;
rule_s_t din_1_20;
rule_s_t din_1_20_r1;
rule_s_t din_1_20_r2;
logic din_valid_1_20;
logic din_valid_1_20_r1;
logic din_valid_1_20_r2;
logic din_ready_1_20;
logic din_almost_full_1_20;
logic [31:0] din_csr_readdata_1_20;
rule_s_t back_data_1_20;
logic    back_valid_1_20;
logic    back_ready_1_20;
logic [RID_WIDTH-1:0] hash_out_1_21;
logic hash_out_valid_filter_1_21;
rule_s_t din_1_21;
rule_s_t din_1_21_r1;
rule_s_t din_1_21_r2;
logic din_valid_1_21;
logic din_valid_1_21_r1;
logic din_valid_1_21_r2;
logic din_ready_1_21;
logic din_almost_full_1_21;
logic [31:0] din_csr_readdata_1_21;
rule_s_t back_data_1_21;
logic    back_valid_1_21;
logic    back_ready_1_21;
logic [RID_WIDTH-1:0] hash_out_1_22;
logic hash_out_valid_filter_1_22;
rule_s_t din_1_22;
rule_s_t din_1_22_r1;
rule_s_t din_1_22_r2;
logic din_valid_1_22;
logic din_valid_1_22_r1;
logic din_valid_1_22_r2;
logic din_ready_1_22;
logic din_almost_full_1_22;
logic [31:0] din_csr_readdata_1_22;
rule_s_t back_data_1_22;
logic    back_valid_1_22;
logic    back_ready_1_22;
logic [RID_WIDTH-1:0] hash_out_1_23;
logic hash_out_valid_filter_1_23;
rule_s_t din_1_23;
rule_s_t din_1_23_r1;
rule_s_t din_1_23_r2;
logic din_valid_1_23;
logic din_valid_1_23_r1;
logic din_valid_1_23_r2;
logic din_ready_1_23;
logic din_almost_full_1_23;
logic [31:0] din_csr_readdata_1_23;
rule_s_t back_data_1_23;
logic    back_valid_1_23;
logic    back_ready_1_23;
logic [RID_WIDTH-1:0] hash_out_1_24;
logic hash_out_valid_filter_1_24;
rule_s_t din_1_24;
rule_s_t din_1_24_r1;
rule_s_t din_1_24_r2;
logic din_valid_1_24;
logic din_valid_1_24_r1;
logic din_valid_1_24_r2;
logic din_ready_1_24;
logic din_almost_full_1_24;
logic [31:0] din_csr_readdata_1_24;
rule_s_t back_data_1_24;
logic    back_valid_1_24;
logic    back_ready_1_24;
logic [RID_WIDTH-1:0] hash_out_1_25;
logic hash_out_valid_filter_1_25;
rule_s_t din_1_25;
rule_s_t din_1_25_r1;
rule_s_t din_1_25_r2;
logic din_valid_1_25;
logic din_valid_1_25_r1;
logic din_valid_1_25_r2;
logic din_ready_1_25;
logic din_almost_full_1_25;
logic [31:0] din_csr_readdata_1_25;
rule_s_t back_data_1_25;
logic    back_valid_1_25;
logic    back_ready_1_25;
logic [RID_WIDTH-1:0] hash_out_1_26;
logic hash_out_valid_filter_1_26;
rule_s_t din_1_26;
rule_s_t din_1_26_r1;
rule_s_t din_1_26_r2;
logic din_valid_1_26;
logic din_valid_1_26_r1;
logic din_valid_1_26_r2;
logic din_ready_1_26;
logic din_almost_full_1_26;
logic [31:0] din_csr_readdata_1_26;
rule_s_t back_data_1_26;
logic    back_valid_1_26;
logic    back_ready_1_26;
logic [RID_WIDTH-1:0] hash_out_1_27;
logic hash_out_valid_filter_1_27;
rule_s_t din_1_27;
rule_s_t din_1_27_r1;
rule_s_t din_1_27_r2;
logic din_valid_1_27;
logic din_valid_1_27_r1;
logic din_valid_1_27_r2;
logic din_ready_1_27;
logic din_almost_full_1_27;
logic [31:0] din_csr_readdata_1_27;
rule_s_t back_data_1_27;
logic    back_valid_1_27;
logic    back_ready_1_27;
logic [RID_WIDTH-1:0] hash_out_1_28;
logic hash_out_valid_filter_1_28;
rule_s_t din_1_28;
rule_s_t din_1_28_r1;
rule_s_t din_1_28_r2;
logic din_valid_1_28;
logic din_valid_1_28_r1;
logic din_valid_1_28_r2;
logic din_ready_1_28;
logic din_almost_full_1_28;
logic [31:0] din_csr_readdata_1_28;
rule_s_t back_data_1_28;
logic    back_valid_1_28;
logic    back_ready_1_28;
logic [RID_WIDTH-1:0] hash_out_1_29;
logic hash_out_valid_filter_1_29;
rule_s_t din_1_29;
rule_s_t din_1_29_r1;
rule_s_t din_1_29_r2;
logic din_valid_1_29;
logic din_valid_1_29_r1;
logic din_valid_1_29_r2;
logic din_ready_1_29;
logic din_almost_full_1_29;
logic [31:0] din_csr_readdata_1_29;
rule_s_t back_data_1_29;
logic    back_valid_1_29;
logic    back_ready_1_29;
logic [RID_WIDTH-1:0] hash_out_1_30;
logic hash_out_valid_filter_1_30;
rule_s_t din_1_30;
rule_s_t din_1_30_r1;
rule_s_t din_1_30_r2;
logic din_valid_1_30;
logic din_valid_1_30_r1;
logic din_valid_1_30_r2;
logic din_ready_1_30;
logic din_almost_full_1_30;
logic [31:0] din_csr_readdata_1_30;
rule_s_t back_data_1_30;
logic    back_valid_1_30;
logic    back_ready_1_30;
logic [RID_WIDTH-1:0] hash_out_1_31;
logic hash_out_valid_filter_1_31;
rule_s_t din_1_31;
rule_s_t din_1_31_r1;
rule_s_t din_1_31_r2;
logic din_valid_1_31;
logic din_valid_1_31_r1;
logic din_valid_1_31_r2;
logic din_ready_1_31;
logic din_almost_full_1_31;
logic [31:0] din_csr_readdata_1_31;
rule_s_t back_data_1_31;
logic    back_valid_1_31;
logic    back_ready_1_31;
logic [RID_WIDTH-1:0] hash_out_2_0;
logic hash_out_valid_filter_2_0;
rule_s_t din_2_0;
rule_s_t din_2_0_r1;
rule_s_t din_2_0_r2;
logic din_valid_2_0;
logic din_valid_2_0_r1;
logic din_valid_2_0_r2;
logic din_ready_2_0;
logic din_almost_full_2_0;
logic [31:0] din_csr_readdata_2_0;
rule_s_t back_data_2_0;
logic    back_valid_2_0;
logic    back_ready_2_0;
logic [RID_WIDTH-1:0] hash_out_2_1;
logic hash_out_valid_filter_2_1;
rule_s_t din_2_1;
rule_s_t din_2_1_r1;
rule_s_t din_2_1_r2;
logic din_valid_2_1;
logic din_valid_2_1_r1;
logic din_valid_2_1_r2;
logic din_ready_2_1;
logic din_almost_full_2_1;
logic [31:0] din_csr_readdata_2_1;
rule_s_t back_data_2_1;
logic    back_valid_2_1;
logic    back_ready_2_1;
logic [RID_WIDTH-1:0] hash_out_2_2;
logic hash_out_valid_filter_2_2;
rule_s_t din_2_2;
rule_s_t din_2_2_r1;
rule_s_t din_2_2_r2;
logic din_valid_2_2;
logic din_valid_2_2_r1;
logic din_valid_2_2_r2;
logic din_ready_2_2;
logic din_almost_full_2_2;
logic [31:0] din_csr_readdata_2_2;
rule_s_t back_data_2_2;
logic    back_valid_2_2;
logic    back_ready_2_2;
logic [RID_WIDTH-1:0] hash_out_2_3;
logic hash_out_valid_filter_2_3;
rule_s_t din_2_3;
rule_s_t din_2_3_r1;
rule_s_t din_2_3_r2;
logic din_valid_2_3;
logic din_valid_2_3_r1;
logic din_valid_2_3_r2;
logic din_ready_2_3;
logic din_almost_full_2_3;
logic [31:0] din_csr_readdata_2_3;
rule_s_t back_data_2_3;
logic    back_valid_2_3;
logic    back_ready_2_3;
logic [RID_WIDTH-1:0] hash_out_2_4;
logic hash_out_valid_filter_2_4;
rule_s_t din_2_4;
rule_s_t din_2_4_r1;
rule_s_t din_2_4_r2;
logic din_valid_2_4;
logic din_valid_2_4_r1;
logic din_valid_2_4_r2;
logic din_ready_2_4;
logic din_almost_full_2_4;
logic [31:0] din_csr_readdata_2_4;
rule_s_t back_data_2_4;
logic    back_valid_2_4;
logic    back_ready_2_4;
logic [RID_WIDTH-1:0] hash_out_2_5;
logic hash_out_valid_filter_2_5;
rule_s_t din_2_5;
rule_s_t din_2_5_r1;
rule_s_t din_2_5_r2;
logic din_valid_2_5;
logic din_valid_2_5_r1;
logic din_valid_2_5_r2;
logic din_ready_2_5;
logic din_almost_full_2_5;
logic [31:0] din_csr_readdata_2_5;
rule_s_t back_data_2_5;
logic    back_valid_2_5;
logic    back_ready_2_5;
logic [RID_WIDTH-1:0] hash_out_2_6;
logic hash_out_valid_filter_2_6;
rule_s_t din_2_6;
rule_s_t din_2_6_r1;
rule_s_t din_2_6_r2;
logic din_valid_2_6;
logic din_valid_2_6_r1;
logic din_valid_2_6_r2;
logic din_ready_2_6;
logic din_almost_full_2_6;
logic [31:0] din_csr_readdata_2_6;
rule_s_t back_data_2_6;
logic    back_valid_2_6;
logic    back_ready_2_6;
logic [RID_WIDTH-1:0] hash_out_2_7;
logic hash_out_valid_filter_2_7;
rule_s_t din_2_7;
rule_s_t din_2_7_r1;
rule_s_t din_2_7_r2;
logic din_valid_2_7;
logic din_valid_2_7_r1;
logic din_valid_2_7_r2;
logic din_ready_2_7;
logic din_almost_full_2_7;
logic [31:0] din_csr_readdata_2_7;
rule_s_t back_data_2_7;
logic    back_valid_2_7;
logic    back_ready_2_7;
logic [RID_WIDTH-1:0] hash_out_2_8;
logic hash_out_valid_filter_2_8;
rule_s_t din_2_8;
rule_s_t din_2_8_r1;
rule_s_t din_2_8_r2;
logic din_valid_2_8;
logic din_valid_2_8_r1;
logic din_valid_2_8_r2;
logic din_ready_2_8;
logic din_almost_full_2_8;
logic [31:0] din_csr_readdata_2_8;
rule_s_t back_data_2_8;
logic    back_valid_2_8;
logic    back_ready_2_8;
logic [RID_WIDTH-1:0] hash_out_2_9;
logic hash_out_valid_filter_2_9;
rule_s_t din_2_9;
rule_s_t din_2_9_r1;
rule_s_t din_2_9_r2;
logic din_valid_2_9;
logic din_valid_2_9_r1;
logic din_valid_2_9_r2;
logic din_ready_2_9;
logic din_almost_full_2_9;
logic [31:0] din_csr_readdata_2_9;
rule_s_t back_data_2_9;
logic    back_valid_2_9;
logic    back_ready_2_9;
logic [RID_WIDTH-1:0] hash_out_2_10;
logic hash_out_valid_filter_2_10;
rule_s_t din_2_10;
rule_s_t din_2_10_r1;
rule_s_t din_2_10_r2;
logic din_valid_2_10;
logic din_valid_2_10_r1;
logic din_valid_2_10_r2;
logic din_ready_2_10;
logic din_almost_full_2_10;
logic [31:0] din_csr_readdata_2_10;
rule_s_t back_data_2_10;
logic    back_valid_2_10;
logic    back_ready_2_10;
logic [RID_WIDTH-1:0] hash_out_2_11;
logic hash_out_valid_filter_2_11;
rule_s_t din_2_11;
rule_s_t din_2_11_r1;
rule_s_t din_2_11_r2;
logic din_valid_2_11;
logic din_valid_2_11_r1;
logic din_valid_2_11_r2;
logic din_ready_2_11;
logic din_almost_full_2_11;
logic [31:0] din_csr_readdata_2_11;
rule_s_t back_data_2_11;
logic    back_valid_2_11;
logic    back_ready_2_11;
logic [RID_WIDTH-1:0] hash_out_2_12;
logic hash_out_valid_filter_2_12;
rule_s_t din_2_12;
rule_s_t din_2_12_r1;
rule_s_t din_2_12_r2;
logic din_valid_2_12;
logic din_valid_2_12_r1;
logic din_valid_2_12_r2;
logic din_ready_2_12;
logic din_almost_full_2_12;
logic [31:0] din_csr_readdata_2_12;
rule_s_t back_data_2_12;
logic    back_valid_2_12;
logic    back_ready_2_12;
logic [RID_WIDTH-1:0] hash_out_2_13;
logic hash_out_valid_filter_2_13;
rule_s_t din_2_13;
rule_s_t din_2_13_r1;
rule_s_t din_2_13_r2;
logic din_valid_2_13;
logic din_valid_2_13_r1;
logic din_valid_2_13_r2;
logic din_ready_2_13;
logic din_almost_full_2_13;
logic [31:0] din_csr_readdata_2_13;
rule_s_t back_data_2_13;
logic    back_valid_2_13;
logic    back_ready_2_13;
logic [RID_WIDTH-1:0] hash_out_2_14;
logic hash_out_valid_filter_2_14;
rule_s_t din_2_14;
rule_s_t din_2_14_r1;
rule_s_t din_2_14_r2;
logic din_valid_2_14;
logic din_valid_2_14_r1;
logic din_valid_2_14_r2;
logic din_ready_2_14;
logic din_almost_full_2_14;
logic [31:0] din_csr_readdata_2_14;
rule_s_t back_data_2_14;
logic    back_valid_2_14;
logic    back_ready_2_14;
logic [RID_WIDTH-1:0] hash_out_2_15;
logic hash_out_valid_filter_2_15;
rule_s_t din_2_15;
rule_s_t din_2_15_r1;
rule_s_t din_2_15_r2;
logic din_valid_2_15;
logic din_valid_2_15_r1;
logic din_valid_2_15_r2;
logic din_ready_2_15;
logic din_almost_full_2_15;
logic [31:0] din_csr_readdata_2_15;
rule_s_t back_data_2_15;
logic    back_valid_2_15;
logic    back_ready_2_15;
logic [RID_WIDTH-1:0] hash_out_2_16;
logic hash_out_valid_filter_2_16;
rule_s_t din_2_16;
rule_s_t din_2_16_r1;
rule_s_t din_2_16_r2;
logic din_valid_2_16;
logic din_valid_2_16_r1;
logic din_valid_2_16_r2;
logic din_ready_2_16;
logic din_almost_full_2_16;
logic [31:0] din_csr_readdata_2_16;
rule_s_t back_data_2_16;
logic    back_valid_2_16;
logic    back_ready_2_16;
logic [RID_WIDTH-1:0] hash_out_2_17;
logic hash_out_valid_filter_2_17;
rule_s_t din_2_17;
rule_s_t din_2_17_r1;
rule_s_t din_2_17_r2;
logic din_valid_2_17;
logic din_valid_2_17_r1;
logic din_valid_2_17_r2;
logic din_ready_2_17;
logic din_almost_full_2_17;
logic [31:0] din_csr_readdata_2_17;
rule_s_t back_data_2_17;
logic    back_valid_2_17;
logic    back_ready_2_17;
logic [RID_WIDTH-1:0] hash_out_2_18;
logic hash_out_valid_filter_2_18;
rule_s_t din_2_18;
rule_s_t din_2_18_r1;
rule_s_t din_2_18_r2;
logic din_valid_2_18;
logic din_valid_2_18_r1;
logic din_valid_2_18_r2;
logic din_ready_2_18;
logic din_almost_full_2_18;
logic [31:0] din_csr_readdata_2_18;
rule_s_t back_data_2_18;
logic    back_valid_2_18;
logic    back_ready_2_18;
logic [RID_WIDTH-1:0] hash_out_2_19;
logic hash_out_valid_filter_2_19;
rule_s_t din_2_19;
rule_s_t din_2_19_r1;
rule_s_t din_2_19_r2;
logic din_valid_2_19;
logic din_valid_2_19_r1;
logic din_valid_2_19_r2;
logic din_ready_2_19;
logic din_almost_full_2_19;
logic [31:0] din_csr_readdata_2_19;
rule_s_t back_data_2_19;
logic    back_valid_2_19;
logic    back_ready_2_19;
logic [RID_WIDTH-1:0] hash_out_2_20;
logic hash_out_valid_filter_2_20;
rule_s_t din_2_20;
rule_s_t din_2_20_r1;
rule_s_t din_2_20_r2;
logic din_valid_2_20;
logic din_valid_2_20_r1;
logic din_valid_2_20_r2;
logic din_ready_2_20;
logic din_almost_full_2_20;
logic [31:0] din_csr_readdata_2_20;
rule_s_t back_data_2_20;
logic    back_valid_2_20;
logic    back_ready_2_20;
logic [RID_WIDTH-1:0] hash_out_2_21;
logic hash_out_valid_filter_2_21;
rule_s_t din_2_21;
rule_s_t din_2_21_r1;
rule_s_t din_2_21_r2;
logic din_valid_2_21;
logic din_valid_2_21_r1;
logic din_valid_2_21_r2;
logic din_ready_2_21;
logic din_almost_full_2_21;
logic [31:0] din_csr_readdata_2_21;
rule_s_t back_data_2_21;
logic    back_valid_2_21;
logic    back_ready_2_21;
logic [RID_WIDTH-1:0] hash_out_2_22;
logic hash_out_valid_filter_2_22;
rule_s_t din_2_22;
rule_s_t din_2_22_r1;
rule_s_t din_2_22_r2;
logic din_valid_2_22;
logic din_valid_2_22_r1;
logic din_valid_2_22_r2;
logic din_ready_2_22;
logic din_almost_full_2_22;
logic [31:0] din_csr_readdata_2_22;
rule_s_t back_data_2_22;
logic    back_valid_2_22;
logic    back_ready_2_22;
logic [RID_WIDTH-1:0] hash_out_2_23;
logic hash_out_valid_filter_2_23;
rule_s_t din_2_23;
rule_s_t din_2_23_r1;
rule_s_t din_2_23_r2;
logic din_valid_2_23;
logic din_valid_2_23_r1;
logic din_valid_2_23_r2;
logic din_ready_2_23;
logic din_almost_full_2_23;
logic [31:0] din_csr_readdata_2_23;
rule_s_t back_data_2_23;
logic    back_valid_2_23;
logic    back_ready_2_23;
logic [RID_WIDTH-1:0] hash_out_2_24;
logic hash_out_valid_filter_2_24;
rule_s_t din_2_24;
rule_s_t din_2_24_r1;
rule_s_t din_2_24_r2;
logic din_valid_2_24;
logic din_valid_2_24_r1;
logic din_valid_2_24_r2;
logic din_ready_2_24;
logic din_almost_full_2_24;
logic [31:0] din_csr_readdata_2_24;
rule_s_t back_data_2_24;
logic    back_valid_2_24;
logic    back_ready_2_24;
logic [RID_WIDTH-1:0] hash_out_2_25;
logic hash_out_valid_filter_2_25;
rule_s_t din_2_25;
rule_s_t din_2_25_r1;
rule_s_t din_2_25_r2;
logic din_valid_2_25;
logic din_valid_2_25_r1;
logic din_valid_2_25_r2;
logic din_ready_2_25;
logic din_almost_full_2_25;
logic [31:0] din_csr_readdata_2_25;
rule_s_t back_data_2_25;
logic    back_valid_2_25;
logic    back_ready_2_25;
logic [RID_WIDTH-1:0] hash_out_2_26;
logic hash_out_valid_filter_2_26;
rule_s_t din_2_26;
rule_s_t din_2_26_r1;
rule_s_t din_2_26_r2;
logic din_valid_2_26;
logic din_valid_2_26_r1;
logic din_valid_2_26_r2;
logic din_ready_2_26;
logic din_almost_full_2_26;
logic [31:0] din_csr_readdata_2_26;
rule_s_t back_data_2_26;
logic    back_valid_2_26;
logic    back_ready_2_26;
logic [RID_WIDTH-1:0] hash_out_2_27;
logic hash_out_valid_filter_2_27;
rule_s_t din_2_27;
rule_s_t din_2_27_r1;
rule_s_t din_2_27_r2;
logic din_valid_2_27;
logic din_valid_2_27_r1;
logic din_valid_2_27_r2;
logic din_ready_2_27;
logic din_almost_full_2_27;
logic [31:0] din_csr_readdata_2_27;
rule_s_t back_data_2_27;
logic    back_valid_2_27;
logic    back_ready_2_27;
logic [RID_WIDTH-1:0] hash_out_2_28;
logic hash_out_valid_filter_2_28;
rule_s_t din_2_28;
rule_s_t din_2_28_r1;
rule_s_t din_2_28_r2;
logic din_valid_2_28;
logic din_valid_2_28_r1;
logic din_valid_2_28_r2;
logic din_ready_2_28;
logic din_almost_full_2_28;
logic [31:0] din_csr_readdata_2_28;
rule_s_t back_data_2_28;
logic    back_valid_2_28;
logic    back_ready_2_28;
logic [RID_WIDTH-1:0] hash_out_2_29;
logic hash_out_valid_filter_2_29;
rule_s_t din_2_29;
rule_s_t din_2_29_r1;
rule_s_t din_2_29_r2;
logic din_valid_2_29;
logic din_valid_2_29_r1;
logic din_valid_2_29_r2;
logic din_ready_2_29;
logic din_almost_full_2_29;
logic [31:0] din_csr_readdata_2_29;
rule_s_t back_data_2_29;
logic    back_valid_2_29;
logic    back_ready_2_29;
logic [RID_WIDTH-1:0] hash_out_2_30;
logic hash_out_valid_filter_2_30;
rule_s_t din_2_30;
rule_s_t din_2_30_r1;
rule_s_t din_2_30_r2;
logic din_valid_2_30;
logic din_valid_2_30_r1;
logic din_valid_2_30_r2;
logic din_ready_2_30;
logic din_almost_full_2_30;
logic [31:0] din_csr_readdata_2_30;
rule_s_t back_data_2_30;
logic    back_valid_2_30;
logic    back_ready_2_30;
logic [RID_WIDTH-1:0] hash_out_2_31;
logic hash_out_valid_filter_2_31;
rule_s_t din_2_31;
rule_s_t din_2_31_r1;
rule_s_t din_2_31_r2;
logic din_valid_2_31;
logic din_valid_2_31_r1;
logic din_valid_2_31_r2;
logic din_ready_2_31;
logic din_almost_full_2_31;
logic [31:0] din_csr_readdata_2_31;
rule_s_t back_data_2_31;
logic    back_valid_2_31;
logic    back_ready_2_31;
logic [RID_WIDTH-1:0] hash_out_3_0;
logic hash_out_valid_filter_3_0;
rule_s_t din_3_0;
rule_s_t din_3_0_r1;
rule_s_t din_3_0_r2;
logic din_valid_3_0;
logic din_valid_3_0_r1;
logic din_valid_3_0_r2;
logic din_ready_3_0;
logic din_almost_full_3_0;
logic [31:0] din_csr_readdata_3_0;
rule_s_t back_data_3_0;
logic    back_valid_3_0;
logic    back_ready_3_0;
logic [RID_WIDTH-1:0] hash_out_3_1;
logic hash_out_valid_filter_3_1;
rule_s_t din_3_1;
rule_s_t din_3_1_r1;
rule_s_t din_3_1_r2;
logic din_valid_3_1;
logic din_valid_3_1_r1;
logic din_valid_3_1_r2;
logic din_ready_3_1;
logic din_almost_full_3_1;
logic [31:0] din_csr_readdata_3_1;
rule_s_t back_data_3_1;
logic    back_valid_3_1;
logic    back_ready_3_1;
logic [RID_WIDTH-1:0] hash_out_3_2;
logic hash_out_valid_filter_3_2;
rule_s_t din_3_2;
rule_s_t din_3_2_r1;
rule_s_t din_3_2_r2;
logic din_valid_3_2;
logic din_valid_3_2_r1;
logic din_valid_3_2_r2;
logic din_ready_3_2;
logic din_almost_full_3_2;
logic [31:0] din_csr_readdata_3_2;
rule_s_t back_data_3_2;
logic    back_valid_3_2;
logic    back_ready_3_2;
logic [RID_WIDTH-1:0] hash_out_3_3;
logic hash_out_valid_filter_3_3;
rule_s_t din_3_3;
rule_s_t din_3_3_r1;
rule_s_t din_3_3_r2;
logic din_valid_3_3;
logic din_valid_3_3_r1;
logic din_valid_3_3_r2;
logic din_ready_3_3;
logic din_almost_full_3_3;
logic [31:0] din_csr_readdata_3_3;
rule_s_t back_data_3_3;
logic    back_valid_3_3;
logic    back_ready_3_3;
logic [RID_WIDTH-1:0] hash_out_3_4;
logic hash_out_valid_filter_3_4;
rule_s_t din_3_4;
rule_s_t din_3_4_r1;
rule_s_t din_3_4_r2;
logic din_valid_3_4;
logic din_valid_3_4_r1;
logic din_valid_3_4_r2;
logic din_ready_3_4;
logic din_almost_full_3_4;
logic [31:0] din_csr_readdata_3_4;
rule_s_t back_data_3_4;
logic    back_valid_3_4;
logic    back_ready_3_4;
logic [RID_WIDTH-1:0] hash_out_3_5;
logic hash_out_valid_filter_3_5;
rule_s_t din_3_5;
rule_s_t din_3_5_r1;
rule_s_t din_3_5_r2;
logic din_valid_3_5;
logic din_valid_3_5_r1;
logic din_valid_3_5_r2;
logic din_ready_3_5;
logic din_almost_full_3_5;
logic [31:0] din_csr_readdata_3_5;
rule_s_t back_data_3_5;
logic    back_valid_3_5;
logic    back_ready_3_5;
logic [RID_WIDTH-1:0] hash_out_3_6;
logic hash_out_valid_filter_3_6;
rule_s_t din_3_6;
rule_s_t din_3_6_r1;
rule_s_t din_3_6_r2;
logic din_valid_3_6;
logic din_valid_3_6_r1;
logic din_valid_3_6_r2;
logic din_ready_3_6;
logic din_almost_full_3_6;
logic [31:0] din_csr_readdata_3_6;
rule_s_t back_data_3_6;
logic    back_valid_3_6;
logic    back_ready_3_6;
logic [RID_WIDTH-1:0] hash_out_3_7;
logic hash_out_valid_filter_3_7;
rule_s_t din_3_7;
rule_s_t din_3_7_r1;
rule_s_t din_3_7_r2;
logic din_valid_3_7;
logic din_valid_3_7_r1;
logic din_valid_3_7_r2;
logic din_ready_3_7;
logic din_almost_full_3_7;
logic [31:0] din_csr_readdata_3_7;
rule_s_t back_data_3_7;
logic    back_valid_3_7;
logic    back_ready_3_7;
logic [RID_WIDTH-1:0] hash_out_3_8;
logic hash_out_valid_filter_3_8;
rule_s_t din_3_8;
rule_s_t din_3_8_r1;
rule_s_t din_3_8_r2;
logic din_valid_3_8;
logic din_valid_3_8_r1;
logic din_valid_3_8_r2;
logic din_ready_3_8;
logic din_almost_full_3_8;
logic [31:0] din_csr_readdata_3_8;
rule_s_t back_data_3_8;
logic    back_valid_3_8;
logic    back_ready_3_8;
logic [RID_WIDTH-1:0] hash_out_3_9;
logic hash_out_valid_filter_3_9;
rule_s_t din_3_9;
rule_s_t din_3_9_r1;
rule_s_t din_3_9_r2;
logic din_valid_3_9;
logic din_valid_3_9_r1;
logic din_valid_3_9_r2;
logic din_ready_3_9;
logic din_almost_full_3_9;
logic [31:0] din_csr_readdata_3_9;
rule_s_t back_data_3_9;
logic    back_valid_3_9;
logic    back_ready_3_9;
logic [RID_WIDTH-1:0] hash_out_3_10;
logic hash_out_valid_filter_3_10;
rule_s_t din_3_10;
rule_s_t din_3_10_r1;
rule_s_t din_3_10_r2;
logic din_valid_3_10;
logic din_valid_3_10_r1;
logic din_valid_3_10_r2;
logic din_ready_3_10;
logic din_almost_full_3_10;
logic [31:0] din_csr_readdata_3_10;
rule_s_t back_data_3_10;
logic    back_valid_3_10;
logic    back_ready_3_10;
logic [RID_WIDTH-1:0] hash_out_3_11;
logic hash_out_valid_filter_3_11;
rule_s_t din_3_11;
rule_s_t din_3_11_r1;
rule_s_t din_3_11_r2;
logic din_valid_3_11;
logic din_valid_3_11_r1;
logic din_valid_3_11_r2;
logic din_ready_3_11;
logic din_almost_full_3_11;
logic [31:0] din_csr_readdata_3_11;
rule_s_t back_data_3_11;
logic    back_valid_3_11;
logic    back_ready_3_11;
logic [RID_WIDTH-1:0] hash_out_3_12;
logic hash_out_valid_filter_3_12;
rule_s_t din_3_12;
rule_s_t din_3_12_r1;
rule_s_t din_3_12_r2;
logic din_valid_3_12;
logic din_valid_3_12_r1;
logic din_valid_3_12_r2;
logic din_ready_3_12;
logic din_almost_full_3_12;
logic [31:0] din_csr_readdata_3_12;
rule_s_t back_data_3_12;
logic    back_valid_3_12;
logic    back_ready_3_12;
logic [RID_WIDTH-1:0] hash_out_3_13;
logic hash_out_valid_filter_3_13;
rule_s_t din_3_13;
rule_s_t din_3_13_r1;
rule_s_t din_3_13_r2;
logic din_valid_3_13;
logic din_valid_3_13_r1;
logic din_valid_3_13_r2;
logic din_ready_3_13;
logic din_almost_full_3_13;
logic [31:0] din_csr_readdata_3_13;
rule_s_t back_data_3_13;
logic    back_valid_3_13;
logic    back_ready_3_13;
logic [RID_WIDTH-1:0] hash_out_3_14;
logic hash_out_valid_filter_3_14;
rule_s_t din_3_14;
rule_s_t din_3_14_r1;
rule_s_t din_3_14_r2;
logic din_valid_3_14;
logic din_valid_3_14_r1;
logic din_valid_3_14_r2;
logic din_ready_3_14;
logic din_almost_full_3_14;
logic [31:0] din_csr_readdata_3_14;
rule_s_t back_data_3_14;
logic    back_valid_3_14;
logic    back_ready_3_14;
logic [RID_WIDTH-1:0] hash_out_3_15;
logic hash_out_valid_filter_3_15;
rule_s_t din_3_15;
rule_s_t din_3_15_r1;
rule_s_t din_3_15_r2;
logic din_valid_3_15;
logic din_valid_3_15_r1;
logic din_valid_3_15_r2;
logic din_ready_3_15;
logic din_almost_full_3_15;
logic [31:0] din_csr_readdata_3_15;
rule_s_t back_data_3_15;
logic    back_valid_3_15;
logic    back_ready_3_15;
logic [RID_WIDTH-1:0] hash_out_3_16;
logic hash_out_valid_filter_3_16;
rule_s_t din_3_16;
rule_s_t din_3_16_r1;
rule_s_t din_3_16_r2;
logic din_valid_3_16;
logic din_valid_3_16_r1;
logic din_valid_3_16_r2;
logic din_ready_3_16;
logic din_almost_full_3_16;
logic [31:0] din_csr_readdata_3_16;
rule_s_t back_data_3_16;
logic    back_valid_3_16;
logic    back_ready_3_16;
logic [RID_WIDTH-1:0] hash_out_3_17;
logic hash_out_valid_filter_3_17;
rule_s_t din_3_17;
rule_s_t din_3_17_r1;
rule_s_t din_3_17_r2;
logic din_valid_3_17;
logic din_valid_3_17_r1;
logic din_valid_3_17_r2;
logic din_ready_3_17;
logic din_almost_full_3_17;
logic [31:0] din_csr_readdata_3_17;
rule_s_t back_data_3_17;
logic    back_valid_3_17;
logic    back_ready_3_17;
logic [RID_WIDTH-1:0] hash_out_3_18;
logic hash_out_valid_filter_3_18;
rule_s_t din_3_18;
rule_s_t din_3_18_r1;
rule_s_t din_3_18_r2;
logic din_valid_3_18;
logic din_valid_3_18_r1;
logic din_valid_3_18_r2;
logic din_ready_3_18;
logic din_almost_full_3_18;
logic [31:0] din_csr_readdata_3_18;
rule_s_t back_data_3_18;
logic    back_valid_3_18;
logic    back_ready_3_18;
logic [RID_WIDTH-1:0] hash_out_3_19;
logic hash_out_valid_filter_3_19;
rule_s_t din_3_19;
rule_s_t din_3_19_r1;
rule_s_t din_3_19_r2;
logic din_valid_3_19;
logic din_valid_3_19_r1;
logic din_valid_3_19_r2;
logic din_ready_3_19;
logic din_almost_full_3_19;
logic [31:0] din_csr_readdata_3_19;
rule_s_t back_data_3_19;
logic    back_valid_3_19;
logic    back_ready_3_19;
logic [RID_WIDTH-1:0] hash_out_3_20;
logic hash_out_valid_filter_3_20;
rule_s_t din_3_20;
rule_s_t din_3_20_r1;
rule_s_t din_3_20_r2;
logic din_valid_3_20;
logic din_valid_3_20_r1;
logic din_valid_3_20_r2;
logic din_ready_3_20;
logic din_almost_full_3_20;
logic [31:0] din_csr_readdata_3_20;
rule_s_t back_data_3_20;
logic    back_valid_3_20;
logic    back_ready_3_20;
logic [RID_WIDTH-1:0] hash_out_3_21;
logic hash_out_valid_filter_3_21;
rule_s_t din_3_21;
rule_s_t din_3_21_r1;
rule_s_t din_3_21_r2;
logic din_valid_3_21;
logic din_valid_3_21_r1;
logic din_valid_3_21_r2;
logic din_ready_3_21;
logic din_almost_full_3_21;
logic [31:0] din_csr_readdata_3_21;
rule_s_t back_data_3_21;
logic    back_valid_3_21;
logic    back_ready_3_21;
logic [RID_WIDTH-1:0] hash_out_3_22;
logic hash_out_valid_filter_3_22;
rule_s_t din_3_22;
rule_s_t din_3_22_r1;
rule_s_t din_3_22_r2;
logic din_valid_3_22;
logic din_valid_3_22_r1;
logic din_valid_3_22_r2;
logic din_ready_3_22;
logic din_almost_full_3_22;
logic [31:0] din_csr_readdata_3_22;
rule_s_t back_data_3_22;
logic    back_valid_3_22;
logic    back_ready_3_22;
logic [RID_WIDTH-1:0] hash_out_3_23;
logic hash_out_valid_filter_3_23;
rule_s_t din_3_23;
rule_s_t din_3_23_r1;
rule_s_t din_3_23_r2;
logic din_valid_3_23;
logic din_valid_3_23_r1;
logic din_valid_3_23_r2;
logic din_ready_3_23;
logic din_almost_full_3_23;
logic [31:0] din_csr_readdata_3_23;
rule_s_t back_data_3_23;
logic    back_valid_3_23;
logic    back_ready_3_23;
logic [RID_WIDTH-1:0] hash_out_3_24;
logic hash_out_valid_filter_3_24;
rule_s_t din_3_24;
rule_s_t din_3_24_r1;
rule_s_t din_3_24_r2;
logic din_valid_3_24;
logic din_valid_3_24_r1;
logic din_valid_3_24_r2;
logic din_ready_3_24;
logic din_almost_full_3_24;
logic [31:0] din_csr_readdata_3_24;
rule_s_t back_data_3_24;
logic    back_valid_3_24;
logic    back_ready_3_24;
logic [RID_WIDTH-1:0] hash_out_3_25;
logic hash_out_valid_filter_3_25;
rule_s_t din_3_25;
rule_s_t din_3_25_r1;
rule_s_t din_3_25_r2;
logic din_valid_3_25;
logic din_valid_3_25_r1;
logic din_valid_3_25_r2;
logic din_ready_3_25;
logic din_almost_full_3_25;
logic [31:0] din_csr_readdata_3_25;
rule_s_t back_data_3_25;
logic    back_valid_3_25;
logic    back_ready_3_25;
logic [RID_WIDTH-1:0] hash_out_3_26;
logic hash_out_valid_filter_3_26;
rule_s_t din_3_26;
rule_s_t din_3_26_r1;
rule_s_t din_3_26_r2;
logic din_valid_3_26;
logic din_valid_3_26_r1;
logic din_valid_3_26_r2;
logic din_ready_3_26;
logic din_almost_full_3_26;
logic [31:0] din_csr_readdata_3_26;
rule_s_t back_data_3_26;
logic    back_valid_3_26;
logic    back_ready_3_26;
logic [RID_WIDTH-1:0] hash_out_3_27;
logic hash_out_valid_filter_3_27;
rule_s_t din_3_27;
rule_s_t din_3_27_r1;
rule_s_t din_3_27_r2;
logic din_valid_3_27;
logic din_valid_3_27_r1;
logic din_valid_3_27_r2;
logic din_ready_3_27;
logic din_almost_full_3_27;
logic [31:0] din_csr_readdata_3_27;
rule_s_t back_data_3_27;
logic    back_valid_3_27;
logic    back_ready_3_27;
logic [RID_WIDTH-1:0] hash_out_3_28;
logic hash_out_valid_filter_3_28;
rule_s_t din_3_28;
rule_s_t din_3_28_r1;
rule_s_t din_3_28_r2;
logic din_valid_3_28;
logic din_valid_3_28_r1;
logic din_valid_3_28_r2;
logic din_ready_3_28;
logic din_almost_full_3_28;
logic [31:0] din_csr_readdata_3_28;
rule_s_t back_data_3_28;
logic    back_valid_3_28;
logic    back_ready_3_28;
logic [RID_WIDTH-1:0] hash_out_3_29;
logic hash_out_valid_filter_3_29;
rule_s_t din_3_29;
rule_s_t din_3_29_r1;
rule_s_t din_3_29_r2;
logic din_valid_3_29;
logic din_valid_3_29_r1;
logic din_valid_3_29_r2;
logic din_ready_3_29;
logic din_almost_full_3_29;
logic [31:0] din_csr_readdata_3_29;
rule_s_t back_data_3_29;
logic    back_valid_3_29;
logic    back_ready_3_29;
logic [RID_WIDTH-1:0] hash_out_3_30;
logic hash_out_valid_filter_3_30;
rule_s_t din_3_30;
rule_s_t din_3_30_r1;
rule_s_t din_3_30_r2;
logic din_valid_3_30;
logic din_valid_3_30_r1;
logic din_valid_3_30_r2;
logic din_ready_3_30;
logic din_almost_full_3_30;
logic [31:0] din_csr_readdata_3_30;
rule_s_t back_data_3_30;
logic    back_valid_3_30;
logic    back_ready_3_30;
logic [RID_WIDTH-1:0] hash_out_3_31;
logic hash_out_valid_filter_3_31;
rule_s_t din_3_31;
rule_s_t din_3_31_r1;
rule_s_t din_3_31_r2;
logic din_valid_3_31;
logic din_valid_3_31_r1;
logic din_valid_3_31_r2;
logic din_ready_3_31;
logic din_almost_full_3_31;
logic [31:0] din_csr_readdata_3_31;
rule_s_t back_data_3_31;
logic    back_valid_3_31;
logic    back_ready_3_31;
logic [RID_WIDTH-1:0] hash_out_4_0;
logic hash_out_valid_filter_4_0;
rule_s_t din_4_0;
rule_s_t din_4_0_r1;
rule_s_t din_4_0_r2;
logic din_valid_4_0;
logic din_valid_4_0_r1;
logic din_valid_4_0_r2;
logic din_ready_4_0;
logic din_almost_full_4_0;
logic [31:0] din_csr_readdata_4_0;
rule_s_t back_data_4_0;
logic    back_valid_4_0;
logic    back_ready_4_0;
logic [RID_WIDTH-1:0] hash_out_4_1;
logic hash_out_valid_filter_4_1;
rule_s_t din_4_1;
rule_s_t din_4_1_r1;
rule_s_t din_4_1_r2;
logic din_valid_4_1;
logic din_valid_4_1_r1;
logic din_valid_4_1_r2;
logic din_ready_4_1;
logic din_almost_full_4_1;
logic [31:0] din_csr_readdata_4_1;
rule_s_t back_data_4_1;
logic    back_valid_4_1;
logic    back_ready_4_1;
logic [RID_WIDTH-1:0] hash_out_4_2;
logic hash_out_valid_filter_4_2;
rule_s_t din_4_2;
rule_s_t din_4_2_r1;
rule_s_t din_4_2_r2;
logic din_valid_4_2;
logic din_valid_4_2_r1;
logic din_valid_4_2_r2;
logic din_ready_4_2;
logic din_almost_full_4_2;
logic [31:0] din_csr_readdata_4_2;
rule_s_t back_data_4_2;
logic    back_valid_4_2;
logic    back_ready_4_2;
logic [RID_WIDTH-1:0] hash_out_4_3;
logic hash_out_valid_filter_4_3;
rule_s_t din_4_3;
rule_s_t din_4_3_r1;
rule_s_t din_4_3_r2;
logic din_valid_4_3;
logic din_valid_4_3_r1;
logic din_valid_4_3_r2;
logic din_ready_4_3;
logic din_almost_full_4_3;
logic [31:0] din_csr_readdata_4_3;
rule_s_t back_data_4_3;
logic    back_valid_4_3;
logic    back_ready_4_3;
logic [RID_WIDTH-1:0] hash_out_4_4;
logic hash_out_valid_filter_4_4;
rule_s_t din_4_4;
rule_s_t din_4_4_r1;
rule_s_t din_4_4_r2;
logic din_valid_4_4;
logic din_valid_4_4_r1;
logic din_valid_4_4_r2;
logic din_ready_4_4;
logic din_almost_full_4_4;
logic [31:0] din_csr_readdata_4_4;
rule_s_t back_data_4_4;
logic    back_valid_4_4;
logic    back_ready_4_4;
logic [RID_WIDTH-1:0] hash_out_4_5;
logic hash_out_valid_filter_4_5;
rule_s_t din_4_5;
rule_s_t din_4_5_r1;
rule_s_t din_4_5_r2;
logic din_valid_4_5;
logic din_valid_4_5_r1;
logic din_valid_4_5_r2;
logic din_ready_4_5;
logic din_almost_full_4_5;
logic [31:0] din_csr_readdata_4_5;
rule_s_t back_data_4_5;
logic    back_valid_4_5;
logic    back_ready_4_5;
logic [RID_WIDTH-1:0] hash_out_4_6;
logic hash_out_valid_filter_4_6;
rule_s_t din_4_6;
rule_s_t din_4_6_r1;
rule_s_t din_4_6_r2;
logic din_valid_4_6;
logic din_valid_4_6_r1;
logic din_valid_4_6_r2;
logic din_ready_4_6;
logic din_almost_full_4_6;
logic [31:0] din_csr_readdata_4_6;
rule_s_t back_data_4_6;
logic    back_valid_4_6;
logic    back_ready_4_6;
logic [RID_WIDTH-1:0] hash_out_4_7;
logic hash_out_valid_filter_4_7;
rule_s_t din_4_7;
rule_s_t din_4_7_r1;
rule_s_t din_4_7_r2;
logic din_valid_4_7;
logic din_valid_4_7_r1;
logic din_valid_4_7_r2;
logic din_ready_4_7;
logic din_almost_full_4_7;
logic [31:0] din_csr_readdata_4_7;
rule_s_t back_data_4_7;
logic    back_valid_4_7;
logic    back_ready_4_7;
logic [RID_WIDTH-1:0] hash_out_4_8;
logic hash_out_valid_filter_4_8;
rule_s_t din_4_8;
rule_s_t din_4_8_r1;
rule_s_t din_4_8_r2;
logic din_valid_4_8;
logic din_valid_4_8_r1;
logic din_valid_4_8_r2;
logic din_ready_4_8;
logic din_almost_full_4_8;
logic [31:0] din_csr_readdata_4_8;
rule_s_t back_data_4_8;
logic    back_valid_4_8;
logic    back_ready_4_8;
logic [RID_WIDTH-1:0] hash_out_4_9;
logic hash_out_valid_filter_4_9;
rule_s_t din_4_9;
rule_s_t din_4_9_r1;
rule_s_t din_4_9_r2;
logic din_valid_4_9;
logic din_valid_4_9_r1;
logic din_valid_4_9_r2;
logic din_ready_4_9;
logic din_almost_full_4_9;
logic [31:0] din_csr_readdata_4_9;
rule_s_t back_data_4_9;
logic    back_valid_4_9;
logic    back_ready_4_9;
logic [RID_WIDTH-1:0] hash_out_4_10;
logic hash_out_valid_filter_4_10;
rule_s_t din_4_10;
rule_s_t din_4_10_r1;
rule_s_t din_4_10_r2;
logic din_valid_4_10;
logic din_valid_4_10_r1;
logic din_valid_4_10_r2;
logic din_ready_4_10;
logic din_almost_full_4_10;
logic [31:0] din_csr_readdata_4_10;
rule_s_t back_data_4_10;
logic    back_valid_4_10;
logic    back_ready_4_10;
logic [RID_WIDTH-1:0] hash_out_4_11;
logic hash_out_valid_filter_4_11;
rule_s_t din_4_11;
rule_s_t din_4_11_r1;
rule_s_t din_4_11_r2;
logic din_valid_4_11;
logic din_valid_4_11_r1;
logic din_valid_4_11_r2;
logic din_ready_4_11;
logic din_almost_full_4_11;
logic [31:0] din_csr_readdata_4_11;
rule_s_t back_data_4_11;
logic    back_valid_4_11;
logic    back_ready_4_11;
logic [RID_WIDTH-1:0] hash_out_4_12;
logic hash_out_valid_filter_4_12;
rule_s_t din_4_12;
rule_s_t din_4_12_r1;
rule_s_t din_4_12_r2;
logic din_valid_4_12;
logic din_valid_4_12_r1;
logic din_valid_4_12_r2;
logic din_ready_4_12;
logic din_almost_full_4_12;
logic [31:0] din_csr_readdata_4_12;
rule_s_t back_data_4_12;
logic    back_valid_4_12;
logic    back_ready_4_12;
logic [RID_WIDTH-1:0] hash_out_4_13;
logic hash_out_valid_filter_4_13;
rule_s_t din_4_13;
rule_s_t din_4_13_r1;
rule_s_t din_4_13_r2;
logic din_valid_4_13;
logic din_valid_4_13_r1;
logic din_valid_4_13_r2;
logic din_ready_4_13;
logic din_almost_full_4_13;
logic [31:0] din_csr_readdata_4_13;
rule_s_t back_data_4_13;
logic    back_valid_4_13;
logic    back_ready_4_13;
logic [RID_WIDTH-1:0] hash_out_4_14;
logic hash_out_valid_filter_4_14;
rule_s_t din_4_14;
rule_s_t din_4_14_r1;
rule_s_t din_4_14_r2;
logic din_valid_4_14;
logic din_valid_4_14_r1;
logic din_valid_4_14_r2;
logic din_ready_4_14;
logic din_almost_full_4_14;
logic [31:0] din_csr_readdata_4_14;
rule_s_t back_data_4_14;
logic    back_valid_4_14;
logic    back_ready_4_14;
logic [RID_WIDTH-1:0] hash_out_4_15;
logic hash_out_valid_filter_4_15;
rule_s_t din_4_15;
rule_s_t din_4_15_r1;
rule_s_t din_4_15_r2;
logic din_valid_4_15;
logic din_valid_4_15_r1;
logic din_valid_4_15_r2;
logic din_ready_4_15;
logic din_almost_full_4_15;
logic [31:0] din_csr_readdata_4_15;
rule_s_t back_data_4_15;
logic    back_valid_4_15;
logic    back_ready_4_15;
logic [RID_WIDTH-1:0] hash_out_4_16;
logic hash_out_valid_filter_4_16;
rule_s_t din_4_16;
rule_s_t din_4_16_r1;
rule_s_t din_4_16_r2;
logic din_valid_4_16;
logic din_valid_4_16_r1;
logic din_valid_4_16_r2;
logic din_ready_4_16;
logic din_almost_full_4_16;
logic [31:0] din_csr_readdata_4_16;
rule_s_t back_data_4_16;
logic    back_valid_4_16;
logic    back_ready_4_16;
logic [RID_WIDTH-1:0] hash_out_4_17;
logic hash_out_valid_filter_4_17;
rule_s_t din_4_17;
rule_s_t din_4_17_r1;
rule_s_t din_4_17_r2;
logic din_valid_4_17;
logic din_valid_4_17_r1;
logic din_valid_4_17_r2;
logic din_ready_4_17;
logic din_almost_full_4_17;
logic [31:0] din_csr_readdata_4_17;
rule_s_t back_data_4_17;
logic    back_valid_4_17;
logic    back_ready_4_17;
logic [RID_WIDTH-1:0] hash_out_4_18;
logic hash_out_valid_filter_4_18;
rule_s_t din_4_18;
rule_s_t din_4_18_r1;
rule_s_t din_4_18_r2;
logic din_valid_4_18;
logic din_valid_4_18_r1;
logic din_valid_4_18_r2;
logic din_ready_4_18;
logic din_almost_full_4_18;
logic [31:0] din_csr_readdata_4_18;
rule_s_t back_data_4_18;
logic    back_valid_4_18;
logic    back_ready_4_18;
logic [RID_WIDTH-1:0] hash_out_4_19;
logic hash_out_valid_filter_4_19;
rule_s_t din_4_19;
rule_s_t din_4_19_r1;
rule_s_t din_4_19_r2;
logic din_valid_4_19;
logic din_valid_4_19_r1;
logic din_valid_4_19_r2;
logic din_ready_4_19;
logic din_almost_full_4_19;
logic [31:0] din_csr_readdata_4_19;
rule_s_t back_data_4_19;
logic    back_valid_4_19;
logic    back_ready_4_19;
logic [RID_WIDTH-1:0] hash_out_4_20;
logic hash_out_valid_filter_4_20;
rule_s_t din_4_20;
rule_s_t din_4_20_r1;
rule_s_t din_4_20_r2;
logic din_valid_4_20;
logic din_valid_4_20_r1;
logic din_valid_4_20_r2;
logic din_ready_4_20;
logic din_almost_full_4_20;
logic [31:0] din_csr_readdata_4_20;
rule_s_t back_data_4_20;
logic    back_valid_4_20;
logic    back_ready_4_20;
logic [RID_WIDTH-1:0] hash_out_4_21;
logic hash_out_valid_filter_4_21;
rule_s_t din_4_21;
rule_s_t din_4_21_r1;
rule_s_t din_4_21_r2;
logic din_valid_4_21;
logic din_valid_4_21_r1;
logic din_valid_4_21_r2;
logic din_ready_4_21;
logic din_almost_full_4_21;
logic [31:0] din_csr_readdata_4_21;
rule_s_t back_data_4_21;
logic    back_valid_4_21;
logic    back_ready_4_21;
logic [RID_WIDTH-1:0] hash_out_4_22;
logic hash_out_valid_filter_4_22;
rule_s_t din_4_22;
rule_s_t din_4_22_r1;
rule_s_t din_4_22_r2;
logic din_valid_4_22;
logic din_valid_4_22_r1;
logic din_valid_4_22_r2;
logic din_ready_4_22;
logic din_almost_full_4_22;
logic [31:0] din_csr_readdata_4_22;
rule_s_t back_data_4_22;
logic    back_valid_4_22;
logic    back_ready_4_22;
logic [RID_WIDTH-1:0] hash_out_4_23;
logic hash_out_valid_filter_4_23;
rule_s_t din_4_23;
rule_s_t din_4_23_r1;
rule_s_t din_4_23_r2;
logic din_valid_4_23;
logic din_valid_4_23_r1;
logic din_valid_4_23_r2;
logic din_ready_4_23;
logic din_almost_full_4_23;
logic [31:0] din_csr_readdata_4_23;
rule_s_t back_data_4_23;
logic    back_valid_4_23;
logic    back_ready_4_23;
logic [RID_WIDTH-1:0] hash_out_4_24;
logic hash_out_valid_filter_4_24;
rule_s_t din_4_24;
rule_s_t din_4_24_r1;
rule_s_t din_4_24_r2;
logic din_valid_4_24;
logic din_valid_4_24_r1;
logic din_valid_4_24_r2;
logic din_ready_4_24;
logic din_almost_full_4_24;
logic [31:0] din_csr_readdata_4_24;
rule_s_t back_data_4_24;
logic    back_valid_4_24;
logic    back_ready_4_24;
logic [RID_WIDTH-1:0] hash_out_4_25;
logic hash_out_valid_filter_4_25;
rule_s_t din_4_25;
rule_s_t din_4_25_r1;
rule_s_t din_4_25_r2;
logic din_valid_4_25;
logic din_valid_4_25_r1;
logic din_valid_4_25_r2;
logic din_ready_4_25;
logic din_almost_full_4_25;
logic [31:0] din_csr_readdata_4_25;
rule_s_t back_data_4_25;
logic    back_valid_4_25;
logic    back_ready_4_25;
logic [RID_WIDTH-1:0] hash_out_4_26;
logic hash_out_valid_filter_4_26;
rule_s_t din_4_26;
rule_s_t din_4_26_r1;
rule_s_t din_4_26_r2;
logic din_valid_4_26;
logic din_valid_4_26_r1;
logic din_valid_4_26_r2;
logic din_ready_4_26;
logic din_almost_full_4_26;
logic [31:0] din_csr_readdata_4_26;
rule_s_t back_data_4_26;
logic    back_valid_4_26;
logic    back_ready_4_26;
logic [RID_WIDTH-1:0] hash_out_4_27;
logic hash_out_valid_filter_4_27;
rule_s_t din_4_27;
rule_s_t din_4_27_r1;
rule_s_t din_4_27_r2;
logic din_valid_4_27;
logic din_valid_4_27_r1;
logic din_valid_4_27_r2;
logic din_ready_4_27;
logic din_almost_full_4_27;
logic [31:0] din_csr_readdata_4_27;
rule_s_t back_data_4_27;
logic    back_valid_4_27;
logic    back_ready_4_27;
logic [RID_WIDTH-1:0] hash_out_4_28;
logic hash_out_valid_filter_4_28;
rule_s_t din_4_28;
rule_s_t din_4_28_r1;
rule_s_t din_4_28_r2;
logic din_valid_4_28;
logic din_valid_4_28_r1;
logic din_valid_4_28_r2;
logic din_ready_4_28;
logic din_almost_full_4_28;
logic [31:0] din_csr_readdata_4_28;
rule_s_t back_data_4_28;
logic    back_valid_4_28;
logic    back_ready_4_28;
logic [RID_WIDTH-1:0] hash_out_4_29;
logic hash_out_valid_filter_4_29;
rule_s_t din_4_29;
rule_s_t din_4_29_r1;
rule_s_t din_4_29_r2;
logic din_valid_4_29;
logic din_valid_4_29_r1;
logic din_valid_4_29_r2;
logic din_ready_4_29;
logic din_almost_full_4_29;
logic [31:0] din_csr_readdata_4_29;
rule_s_t back_data_4_29;
logic    back_valid_4_29;
logic    back_ready_4_29;
logic [RID_WIDTH-1:0] hash_out_4_30;
logic hash_out_valid_filter_4_30;
rule_s_t din_4_30;
rule_s_t din_4_30_r1;
rule_s_t din_4_30_r2;
logic din_valid_4_30;
logic din_valid_4_30_r1;
logic din_valid_4_30_r2;
logic din_ready_4_30;
logic din_almost_full_4_30;
logic [31:0] din_csr_readdata_4_30;
rule_s_t back_data_4_30;
logic    back_valid_4_30;
logic    back_ready_4_30;
logic [RID_WIDTH-1:0] hash_out_4_31;
logic hash_out_valid_filter_4_31;
rule_s_t din_4_31;
rule_s_t din_4_31_r1;
rule_s_t din_4_31_r2;
logic din_valid_4_31;
logic din_valid_4_31_r1;
logic din_valid_4_31_r2;
logic din_ready_4_31;
logic din_almost_full_4_31;
logic [31:0] din_csr_readdata_4_31;
rule_s_t back_data_4_31;
logic    back_valid_4_31;
logic    back_ready_4_31;
logic [RID_WIDTH-1:0] hash_out_5_0;
logic hash_out_valid_filter_5_0;
rule_s_t din_5_0;
rule_s_t din_5_0_r1;
rule_s_t din_5_0_r2;
logic din_valid_5_0;
logic din_valid_5_0_r1;
logic din_valid_5_0_r2;
logic din_ready_5_0;
logic din_almost_full_5_0;
logic [31:0] din_csr_readdata_5_0;
rule_s_t back_data_5_0;
logic    back_valid_5_0;
logic    back_ready_5_0;
logic [RID_WIDTH-1:0] hash_out_5_1;
logic hash_out_valid_filter_5_1;
rule_s_t din_5_1;
rule_s_t din_5_1_r1;
rule_s_t din_5_1_r2;
logic din_valid_5_1;
logic din_valid_5_1_r1;
logic din_valid_5_1_r2;
logic din_ready_5_1;
logic din_almost_full_5_1;
logic [31:0] din_csr_readdata_5_1;
rule_s_t back_data_5_1;
logic    back_valid_5_1;
logic    back_ready_5_1;
logic [RID_WIDTH-1:0] hash_out_5_2;
logic hash_out_valid_filter_5_2;
rule_s_t din_5_2;
rule_s_t din_5_2_r1;
rule_s_t din_5_2_r2;
logic din_valid_5_2;
logic din_valid_5_2_r1;
logic din_valid_5_2_r2;
logic din_ready_5_2;
logic din_almost_full_5_2;
logic [31:0] din_csr_readdata_5_2;
rule_s_t back_data_5_2;
logic    back_valid_5_2;
logic    back_ready_5_2;
logic [RID_WIDTH-1:0] hash_out_5_3;
logic hash_out_valid_filter_5_3;
rule_s_t din_5_3;
rule_s_t din_5_3_r1;
rule_s_t din_5_3_r2;
logic din_valid_5_3;
logic din_valid_5_3_r1;
logic din_valid_5_3_r2;
logic din_ready_5_3;
logic din_almost_full_5_3;
logic [31:0] din_csr_readdata_5_3;
rule_s_t back_data_5_3;
logic    back_valid_5_3;
logic    back_ready_5_3;
logic [RID_WIDTH-1:0] hash_out_5_4;
logic hash_out_valid_filter_5_4;
rule_s_t din_5_4;
rule_s_t din_5_4_r1;
rule_s_t din_5_4_r2;
logic din_valid_5_4;
logic din_valid_5_4_r1;
logic din_valid_5_4_r2;
logic din_ready_5_4;
logic din_almost_full_5_4;
logic [31:0] din_csr_readdata_5_4;
rule_s_t back_data_5_4;
logic    back_valid_5_4;
logic    back_ready_5_4;
logic [RID_WIDTH-1:0] hash_out_5_5;
logic hash_out_valid_filter_5_5;
rule_s_t din_5_5;
rule_s_t din_5_5_r1;
rule_s_t din_5_5_r2;
logic din_valid_5_5;
logic din_valid_5_5_r1;
logic din_valid_5_5_r2;
logic din_ready_5_5;
logic din_almost_full_5_5;
logic [31:0] din_csr_readdata_5_5;
rule_s_t back_data_5_5;
logic    back_valid_5_5;
logic    back_ready_5_5;
logic [RID_WIDTH-1:0] hash_out_5_6;
logic hash_out_valid_filter_5_6;
rule_s_t din_5_6;
rule_s_t din_5_6_r1;
rule_s_t din_5_6_r2;
logic din_valid_5_6;
logic din_valid_5_6_r1;
logic din_valid_5_6_r2;
logic din_ready_5_6;
logic din_almost_full_5_6;
logic [31:0] din_csr_readdata_5_6;
rule_s_t back_data_5_6;
logic    back_valid_5_6;
logic    back_ready_5_6;
logic [RID_WIDTH-1:0] hash_out_5_7;
logic hash_out_valid_filter_5_7;
rule_s_t din_5_7;
rule_s_t din_5_7_r1;
rule_s_t din_5_7_r2;
logic din_valid_5_7;
logic din_valid_5_7_r1;
logic din_valid_5_7_r2;
logic din_ready_5_7;
logic din_almost_full_5_7;
logic [31:0] din_csr_readdata_5_7;
rule_s_t back_data_5_7;
logic    back_valid_5_7;
logic    back_ready_5_7;
logic [RID_WIDTH-1:0] hash_out_5_8;
logic hash_out_valid_filter_5_8;
rule_s_t din_5_8;
rule_s_t din_5_8_r1;
rule_s_t din_5_8_r2;
logic din_valid_5_8;
logic din_valid_5_8_r1;
logic din_valid_5_8_r2;
logic din_ready_5_8;
logic din_almost_full_5_8;
logic [31:0] din_csr_readdata_5_8;
rule_s_t back_data_5_8;
logic    back_valid_5_8;
logic    back_ready_5_8;
logic [RID_WIDTH-1:0] hash_out_5_9;
logic hash_out_valid_filter_5_9;
rule_s_t din_5_9;
rule_s_t din_5_9_r1;
rule_s_t din_5_9_r2;
logic din_valid_5_9;
logic din_valid_5_9_r1;
logic din_valid_5_9_r2;
logic din_ready_5_9;
logic din_almost_full_5_9;
logic [31:0] din_csr_readdata_5_9;
rule_s_t back_data_5_9;
logic    back_valid_5_9;
logic    back_ready_5_9;
logic [RID_WIDTH-1:0] hash_out_5_10;
logic hash_out_valid_filter_5_10;
rule_s_t din_5_10;
rule_s_t din_5_10_r1;
rule_s_t din_5_10_r2;
logic din_valid_5_10;
logic din_valid_5_10_r1;
logic din_valid_5_10_r2;
logic din_ready_5_10;
logic din_almost_full_5_10;
logic [31:0] din_csr_readdata_5_10;
rule_s_t back_data_5_10;
logic    back_valid_5_10;
logic    back_ready_5_10;
logic [RID_WIDTH-1:0] hash_out_5_11;
logic hash_out_valid_filter_5_11;
rule_s_t din_5_11;
rule_s_t din_5_11_r1;
rule_s_t din_5_11_r2;
logic din_valid_5_11;
logic din_valid_5_11_r1;
logic din_valid_5_11_r2;
logic din_ready_5_11;
logic din_almost_full_5_11;
logic [31:0] din_csr_readdata_5_11;
rule_s_t back_data_5_11;
logic    back_valid_5_11;
logic    back_ready_5_11;
logic [RID_WIDTH-1:0] hash_out_5_12;
logic hash_out_valid_filter_5_12;
rule_s_t din_5_12;
rule_s_t din_5_12_r1;
rule_s_t din_5_12_r2;
logic din_valid_5_12;
logic din_valid_5_12_r1;
logic din_valid_5_12_r2;
logic din_ready_5_12;
logic din_almost_full_5_12;
logic [31:0] din_csr_readdata_5_12;
rule_s_t back_data_5_12;
logic    back_valid_5_12;
logic    back_ready_5_12;
logic [RID_WIDTH-1:0] hash_out_5_13;
logic hash_out_valid_filter_5_13;
rule_s_t din_5_13;
rule_s_t din_5_13_r1;
rule_s_t din_5_13_r2;
logic din_valid_5_13;
logic din_valid_5_13_r1;
logic din_valid_5_13_r2;
logic din_ready_5_13;
logic din_almost_full_5_13;
logic [31:0] din_csr_readdata_5_13;
rule_s_t back_data_5_13;
logic    back_valid_5_13;
logic    back_ready_5_13;
logic [RID_WIDTH-1:0] hash_out_5_14;
logic hash_out_valid_filter_5_14;
rule_s_t din_5_14;
rule_s_t din_5_14_r1;
rule_s_t din_5_14_r2;
logic din_valid_5_14;
logic din_valid_5_14_r1;
logic din_valid_5_14_r2;
logic din_ready_5_14;
logic din_almost_full_5_14;
logic [31:0] din_csr_readdata_5_14;
rule_s_t back_data_5_14;
logic    back_valid_5_14;
logic    back_ready_5_14;
logic [RID_WIDTH-1:0] hash_out_5_15;
logic hash_out_valid_filter_5_15;
rule_s_t din_5_15;
rule_s_t din_5_15_r1;
rule_s_t din_5_15_r2;
logic din_valid_5_15;
logic din_valid_5_15_r1;
logic din_valid_5_15_r2;
logic din_ready_5_15;
logic din_almost_full_5_15;
logic [31:0] din_csr_readdata_5_15;
rule_s_t back_data_5_15;
logic    back_valid_5_15;
logic    back_ready_5_15;
logic [RID_WIDTH-1:0] hash_out_5_16;
logic hash_out_valid_filter_5_16;
rule_s_t din_5_16;
rule_s_t din_5_16_r1;
rule_s_t din_5_16_r2;
logic din_valid_5_16;
logic din_valid_5_16_r1;
logic din_valid_5_16_r2;
logic din_ready_5_16;
logic din_almost_full_5_16;
logic [31:0] din_csr_readdata_5_16;
rule_s_t back_data_5_16;
logic    back_valid_5_16;
logic    back_ready_5_16;
logic [RID_WIDTH-1:0] hash_out_5_17;
logic hash_out_valid_filter_5_17;
rule_s_t din_5_17;
rule_s_t din_5_17_r1;
rule_s_t din_5_17_r2;
logic din_valid_5_17;
logic din_valid_5_17_r1;
logic din_valid_5_17_r2;
logic din_ready_5_17;
logic din_almost_full_5_17;
logic [31:0] din_csr_readdata_5_17;
rule_s_t back_data_5_17;
logic    back_valid_5_17;
logic    back_ready_5_17;
logic [RID_WIDTH-1:0] hash_out_5_18;
logic hash_out_valid_filter_5_18;
rule_s_t din_5_18;
rule_s_t din_5_18_r1;
rule_s_t din_5_18_r2;
logic din_valid_5_18;
logic din_valid_5_18_r1;
logic din_valid_5_18_r2;
logic din_ready_5_18;
logic din_almost_full_5_18;
logic [31:0] din_csr_readdata_5_18;
rule_s_t back_data_5_18;
logic    back_valid_5_18;
logic    back_ready_5_18;
logic [RID_WIDTH-1:0] hash_out_5_19;
logic hash_out_valid_filter_5_19;
rule_s_t din_5_19;
rule_s_t din_5_19_r1;
rule_s_t din_5_19_r2;
logic din_valid_5_19;
logic din_valid_5_19_r1;
logic din_valid_5_19_r2;
logic din_ready_5_19;
logic din_almost_full_5_19;
logic [31:0] din_csr_readdata_5_19;
rule_s_t back_data_5_19;
logic    back_valid_5_19;
logic    back_ready_5_19;
logic [RID_WIDTH-1:0] hash_out_5_20;
logic hash_out_valid_filter_5_20;
rule_s_t din_5_20;
rule_s_t din_5_20_r1;
rule_s_t din_5_20_r2;
logic din_valid_5_20;
logic din_valid_5_20_r1;
logic din_valid_5_20_r2;
logic din_ready_5_20;
logic din_almost_full_5_20;
logic [31:0] din_csr_readdata_5_20;
rule_s_t back_data_5_20;
logic    back_valid_5_20;
logic    back_ready_5_20;
logic [RID_WIDTH-1:0] hash_out_5_21;
logic hash_out_valid_filter_5_21;
rule_s_t din_5_21;
rule_s_t din_5_21_r1;
rule_s_t din_5_21_r2;
logic din_valid_5_21;
logic din_valid_5_21_r1;
logic din_valid_5_21_r2;
logic din_ready_5_21;
logic din_almost_full_5_21;
logic [31:0] din_csr_readdata_5_21;
rule_s_t back_data_5_21;
logic    back_valid_5_21;
logic    back_ready_5_21;
logic [RID_WIDTH-1:0] hash_out_5_22;
logic hash_out_valid_filter_5_22;
rule_s_t din_5_22;
rule_s_t din_5_22_r1;
rule_s_t din_5_22_r2;
logic din_valid_5_22;
logic din_valid_5_22_r1;
logic din_valid_5_22_r2;
logic din_ready_5_22;
logic din_almost_full_5_22;
logic [31:0] din_csr_readdata_5_22;
rule_s_t back_data_5_22;
logic    back_valid_5_22;
logic    back_ready_5_22;
logic [RID_WIDTH-1:0] hash_out_5_23;
logic hash_out_valid_filter_5_23;
rule_s_t din_5_23;
rule_s_t din_5_23_r1;
rule_s_t din_5_23_r2;
logic din_valid_5_23;
logic din_valid_5_23_r1;
logic din_valid_5_23_r2;
logic din_ready_5_23;
logic din_almost_full_5_23;
logic [31:0] din_csr_readdata_5_23;
rule_s_t back_data_5_23;
logic    back_valid_5_23;
logic    back_ready_5_23;
logic [RID_WIDTH-1:0] hash_out_5_24;
logic hash_out_valid_filter_5_24;
rule_s_t din_5_24;
rule_s_t din_5_24_r1;
rule_s_t din_5_24_r2;
logic din_valid_5_24;
logic din_valid_5_24_r1;
logic din_valid_5_24_r2;
logic din_ready_5_24;
logic din_almost_full_5_24;
logic [31:0] din_csr_readdata_5_24;
rule_s_t back_data_5_24;
logic    back_valid_5_24;
logic    back_ready_5_24;
logic [RID_WIDTH-1:0] hash_out_5_25;
logic hash_out_valid_filter_5_25;
rule_s_t din_5_25;
rule_s_t din_5_25_r1;
rule_s_t din_5_25_r2;
logic din_valid_5_25;
logic din_valid_5_25_r1;
logic din_valid_5_25_r2;
logic din_ready_5_25;
logic din_almost_full_5_25;
logic [31:0] din_csr_readdata_5_25;
rule_s_t back_data_5_25;
logic    back_valid_5_25;
logic    back_ready_5_25;
logic [RID_WIDTH-1:0] hash_out_5_26;
logic hash_out_valid_filter_5_26;
rule_s_t din_5_26;
rule_s_t din_5_26_r1;
rule_s_t din_5_26_r2;
logic din_valid_5_26;
logic din_valid_5_26_r1;
logic din_valid_5_26_r2;
logic din_ready_5_26;
logic din_almost_full_5_26;
logic [31:0] din_csr_readdata_5_26;
rule_s_t back_data_5_26;
logic    back_valid_5_26;
logic    back_ready_5_26;
logic [RID_WIDTH-1:0] hash_out_5_27;
logic hash_out_valid_filter_5_27;
rule_s_t din_5_27;
rule_s_t din_5_27_r1;
rule_s_t din_5_27_r2;
logic din_valid_5_27;
logic din_valid_5_27_r1;
logic din_valid_5_27_r2;
logic din_ready_5_27;
logic din_almost_full_5_27;
logic [31:0] din_csr_readdata_5_27;
rule_s_t back_data_5_27;
logic    back_valid_5_27;
logic    back_ready_5_27;
logic [RID_WIDTH-1:0] hash_out_5_28;
logic hash_out_valid_filter_5_28;
rule_s_t din_5_28;
rule_s_t din_5_28_r1;
rule_s_t din_5_28_r2;
logic din_valid_5_28;
logic din_valid_5_28_r1;
logic din_valid_5_28_r2;
logic din_ready_5_28;
logic din_almost_full_5_28;
logic [31:0] din_csr_readdata_5_28;
rule_s_t back_data_5_28;
logic    back_valid_5_28;
logic    back_ready_5_28;
logic [RID_WIDTH-1:0] hash_out_5_29;
logic hash_out_valid_filter_5_29;
rule_s_t din_5_29;
rule_s_t din_5_29_r1;
rule_s_t din_5_29_r2;
logic din_valid_5_29;
logic din_valid_5_29_r1;
logic din_valid_5_29_r2;
logic din_ready_5_29;
logic din_almost_full_5_29;
logic [31:0] din_csr_readdata_5_29;
rule_s_t back_data_5_29;
logic    back_valid_5_29;
logic    back_ready_5_29;
logic [RID_WIDTH-1:0] hash_out_5_30;
logic hash_out_valid_filter_5_30;
rule_s_t din_5_30;
rule_s_t din_5_30_r1;
rule_s_t din_5_30_r2;
logic din_valid_5_30;
logic din_valid_5_30_r1;
logic din_valid_5_30_r2;
logic din_ready_5_30;
logic din_almost_full_5_30;
logic [31:0] din_csr_readdata_5_30;
rule_s_t back_data_5_30;
logic    back_valid_5_30;
logic    back_ready_5_30;
logic [RID_WIDTH-1:0] hash_out_5_31;
logic hash_out_valid_filter_5_31;
rule_s_t din_5_31;
rule_s_t din_5_31_r1;
rule_s_t din_5_31_r2;
logic din_valid_5_31;
logic din_valid_5_31_r1;
logic din_valid_5_31_r2;
logic din_ready_5_31;
logic din_almost_full_5_31;
logic [31:0] din_csr_readdata_5_31;
rule_s_t back_data_5_31;
logic    back_valid_5_31;
logic    back_ready_5_31;
logic [RID_WIDTH-1:0] hash_out_6_0;
logic hash_out_valid_filter_6_0;
rule_s_t din_6_0;
rule_s_t din_6_0_r1;
rule_s_t din_6_0_r2;
logic din_valid_6_0;
logic din_valid_6_0_r1;
logic din_valid_6_0_r2;
logic din_ready_6_0;
logic din_almost_full_6_0;
logic [31:0] din_csr_readdata_6_0;
rule_s_t back_data_6_0;
logic    back_valid_6_0;
logic    back_ready_6_0;
logic [RID_WIDTH-1:0] hash_out_6_1;
logic hash_out_valid_filter_6_1;
rule_s_t din_6_1;
rule_s_t din_6_1_r1;
rule_s_t din_6_1_r2;
logic din_valid_6_1;
logic din_valid_6_1_r1;
logic din_valid_6_1_r2;
logic din_ready_6_1;
logic din_almost_full_6_1;
logic [31:0] din_csr_readdata_6_1;
rule_s_t back_data_6_1;
logic    back_valid_6_1;
logic    back_ready_6_1;
logic [RID_WIDTH-1:0] hash_out_6_2;
logic hash_out_valid_filter_6_2;
rule_s_t din_6_2;
rule_s_t din_6_2_r1;
rule_s_t din_6_2_r2;
logic din_valid_6_2;
logic din_valid_6_2_r1;
logic din_valid_6_2_r2;
logic din_ready_6_2;
logic din_almost_full_6_2;
logic [31:0] din_csr_readdata_6_2;
rule_s_t back_data_6_2;
logic    back_valid_6_2;
logic    back_ready_6_2;
logic [RID_WIDTH-1:0] hash_out_6_3;
logic hash_out_valid_filter_6_3;
rule_s_t din_6_3;
rule_s_t din_6_3_r1;
rule_s_t din_6_3_r2;
logic din_valid_6_3;
logic din_valid_6_3_r1;
logic din_valid_6_3_r2;
logic din_ready_6_3;
logic din_almost_full_6_3;
logic [31:0] din_csr_readdata_6_3;
rule_s_t back_data_6_3;
logic    back_valid_6_3;
logic    back_ready_6_3;
logic [RID_WIDTH-1:0] hash_out_6_4;
logic hash_out_valid_filter_6_4;
rule_s_t din_6_4;
rule_s_t din_6_4_r1;
rule_s_t din_6_4_r2;
logic din_valid_6_4;
logic din_valid_6_4_r1;
logic din_valid_6_4_r2;
logic din_ready_6_4;
logic din_almost_full_6_4;
logic [31:0] din_csr_readdata_6_4;
rule_s_t back_data_6_4;
logic    back_valid_6_4;
logic    back_ready_6_4;
logic [RID_WIDTH-1:0] hash_out_6_5;
logic hash_out_valid_filter_6_5;
rule_s_t din_6_5;
rule_s_t din_6_5_r1;
rule_s_t din_6_5_r2;
logic din_valid_6_5;
logic din_valid_6_5_r1;
logic din_valid_6_5_r2;
logic din_ready_6_5;
logic din_almost_full_6_5;
logic [31:0] din_csr_readdata_6_5;
rule_s_t back_data_6_5;
logic    back_valid_6_5;
logic    back_ready_6_5;
logic [RID_WIDTH-1:0] hash_out_6_6;
logic hash_out_valid_filter_6_6;
rule_s_t din_6_6;
rule_s_t din_6_6_r1;
rule_s_t din_6_6_r2;
logic din_valid_6_6;
logic din_valid_6_6_r1;
logic din_valid_6_6_r2;
logic din_ready_6_6;
logic din_almost_full_6_6;
logic [31:0] din_csr_readdata_6_6;
rule_s_t back_data_6_6;
logic    back_valid_6_6;
logic    back_ready_6_6;
logic [RID_WIDTH-1:0] hash_out_6_7;
logic hash_out_valid_filter_6_7;
rule_s_t din_6_7;
rule_s_t din_6_7_r1;
rule_s_t din_6_7_r2;
logic din_valid_6_7;
logic din_valid_6_7_r1;
logic din_valid_6_7_r2;
logic din_ready_6_7;
logic din_almost_full_6_7;
logic [31:0] din_csr_readdata_6_7;
rule_s_t back_data_6_7;
logic    back_valid_6_7;
logic    back_ready_6_7;
logic [RID_WIDTH-1:0] hash_out_6_8;
logic hash_out_valid_filter_6_8;
rule_s_t din_6_8;
rule_s_t din_6_8_r1;
rule_s_t din_6_8_r2;
logic din_valid_6_8;
logic din_valid_6_8_r1;
logic din_valid_6_8_r2;
logic din_ready_6_8;
logic din_almost_full_6_8;
logic [31:0] din_csr_readdata_6_8;
rule_s_t back_data_6_8;
logic    back_valid_6_8;
logic    back_ready_6_8;
logic [RID_WIDTH-1:0] hash_out_6_9;
logic hash_out_valid_filter_6_9;
rule_s_t din_6_9;
rule_s_t din_6_9_r1;
rule_s_t din_6_9_r2;
logic din_valid_6_9;
logic din_valid_6_9_r1;
logic din_valid_6_9_r2;
logic din_ready_6_9;
logic din_almost_full_6_9;
logic [31:0] din_csr_readdata_6_9;
rule_s_t back_data_6_9;
logic    back_valid_6_9;
logic    back_ready_6_9;
logic [RID_WIDTH-1:0] hash_out_6_10;
logic hash_out_valid_filter_6_10;
rule_s_t din_6_10;
rule_s_t din_6_10_r1;
rule_s_t din_6_10_r2;
logic din_valid_6_10;
logic din_valid_6_10_r1;
logic din_valid_6_10_r2;
logic din_ready_6_10;
logic din_almost_full_6_10;
logic [31:0] din_csr_readdata_6_10;
rule_s_t back_data_6_10;
logic    back_valid_6_10;
logic    back_ready_6_10;
logic [RID_WIDTH-1:0] hash_out_6_11;
logic hash_out_valid_filter_6_11;
rule_s_t din_6_11;
rule_s_t din_6_11_r1;
rule_s_t din_6_11_r2;
logic din_valid_6_11;
logic din_valid_6_11_r1;
logic din_valid_6_11_r2;
logic din_ready_6_11;
logic din_almost_full_6_11;
logic [31:0] din_csr_readdata_6_11;
rule_s_t back_data_6_11;
logic    back_valid_6_11;
logic    back_ready_6_11;
logic [RID_WIDTH-1:0] hash_out_6_12;
logic hash_out_valid_filter_6_12;
rule_s_t din_6_12;
rule_s_t din_6_12_r1;
rule_s_t din_6_12_r2;
logic din_valid_6_12;
logic din_valid_6_12_r1;
logic din_valid_6_12_r2;
logic din_ready_6_12;
logic din_almost_full_6_12;
logic [31:0] din_csr_readdata_6_12;
rule_s_t back_data_6_12;
logic    back_valid_6_12;
logic    back_ready_6_12;
logic [RID_WIDTH-1:0] hash_out_6_13;
logic hash_out_valid_filter_6_13;
rule_s_t din_6_13;
rule_s_t din_6_13_r1;
rule_s_t din_6_13_r2;
logic din_valid_6_13;
logic din_valid_6_13_r1;
logic din_valid_6_13_r2;
logic din_ready_6_13;
logic din_almost_full_6_13;
logic [31:0] din_csr_readdata_6_13;
rule_s_t back_data_6_13;
logic    back_valid_6_13;
logic    back_ready_6_13;
logic [RID_WIDTH-1:0] hash_out_6_14;
logic hash_out_valid_filter_6_14;
rule_s_t din_6_14;
rule_s_t din_6_14_r1;
rule_s_t din_6_14_r2;
logic din_valid_6_14;
logic din_valid_6_14_r1;
logic din_valid_6_14_r2;
logic din_ready_6_14;
logic din_almost_full_6_14;
logic [31:0] din_csr_readdata_6_14;
rule_s_t back_data_6_14;
logic    back_valid_6_14;
logic    back_ready_6_14;
logic [RID_WIDTH-1:0] hash_out_6_15;
logic hash_out_valid_filter_6_15;
rule_s_t din_6_15;
rule_s_t din_6_15_r1;
rule_s_t din_6_15_r2;
logic din_valid_6_15;
logic din_valid_6_15_r1;
logic din_valid_6_15_r2;
logic din_ready_6_15;
logic din_almost_full_6_15;
logic [31:0] din_csr_readdata_6_15;
rule_s_t back_data_6_15;
logic    back_valid_6_15;
logic    back_ready_6_15;
logic [RID_WIDTH-1:0] hash_out_6_16;
logic hash_out_valid_filter_6_16;
rule_s_t din_6_16;
rule_s_t din_6_16_r1;
rule_s_t din_6_16_r2;
logic din_valid_6_16;
logic din_valid_6_16_r1;
logic din_valid_6_16_r2;
logic din_ready_6_16;
logic din_almost_full_6_16;
logic [31:0] din_csr_readdata_6_16;
rule_s_t back_data_6_16;
logic    back_valid_6_16;
logic    back_ready_6_16;
logic [RID_WIDTH-1:0] hash_out_6_17;
logic hash_out_valid_filter_6_17;
rule_s_t din_6_17;
rule_s_t din_6_17_r1;
rule_s_t din_6_17_r2;
logic din_valid_6_17;
logic din_valid_6_17_r1;
logic din_valid_6_17_r2;
logic din_ready_6_17;
logic din_almost_full_6_17;
logic [31:0] din_csr_readdata_6_17;
rule_s_t back_data_6_17;
logic    back_valid_6_17;
logic    back_ready_6_17;
logic [RID_WIDTH-1:0] hash_out_6_18;
logic hash_out_valid_filter_6_18;
rule_s_t din_6_18;
rule_s_t din_6_18_r1;
rule_s_t din_6_18_r2;
logic din_valid_6_18;
logic din_valid_6_18_r1;
logic din_valid_6_18_r2;
logic din_ready_6_18;
logic din_almost_full_6_18;
logic [31:0] din_csr_readdata_6_18;
rule_s_t back_data_6_18;
logic    back_valid_6_18;
logic    back_ready_6_18;
logic [RID_WIDTH-1:0] hash_out_6_19;
logic hash_out_valid_filter_6_19;
rule_s_t din_6_19;
rule_s_t din_6_19_r1;
rule_s_t din_6_19_r2;
logic din_valid_6_19;
logic din_valid_6_19_r1;
logic din_valid_6_19_r2;
logic din_ready_6_19;
logic din_almost_full_6_19;
logic [31:0] din_csr_readdata_6_19;
rule_s_t back_data_6_19;
logic    back_valid_6_19;
logic    back_ready_6_19;
logic [RID_WIDTH-1:0] hash_out_6_20;
logic hash_out_valid_filter_6_20;
rule_s_t din_6_20;
rule_s_t din_6_20_r1;
rule_s_t din_6_20_r2;
logic din_valid_6_20;
logic din_valid_6_20_r1;
logic din_valid_6_20_r2;
logic din_ready_6_20;
logic din_almost_full_6_20;
logic [31:0] din_csr_readdata_6_20;
rule_s_t back_data_6_20;
logic    back_valid_6_20;
logic    back_ready_6_20;
logic [RID_WIDTH-1:0] hash_out_6_21;
logic hash_out_valid_filter_6_21;
rule_s_t din_6_21;
rule_s_t din_6_21_r1;
rule_s_t din_6_21_r2;
logic din_valid_6_21;
logic din_valid_6_21_r1;
logic din_valid_6_21_r2;
logic din_ready_6_21;
logic din_almost_full_6_21;
logic [31:0] din_csr_readdata_6_21;
rule_s_t back_data_6_21;
logic    back_valid_6_21;
logic    back_ready_6_21;
logic [RID_WIDTH-1:0] hash_out_6_22;
logic hash_out_valid_filter_6_22;
rule_s_t din_6_22;
rule_s_t din_6_22_r1;
rule_s_t din_6_22_r2;
logic din_valid_6_22;
logic din_valid_6_22_r1;
logic din_valid_6_22_r2;
logic din_ready_6_22;
logic din_almost_full_6_22;
logic [31:0] din_csr_readdata_6_22;
rule_s_t back_data_6_22;
logic    back_valid_6_22;
logic    back_ready_6_22;
logic [RID_WIDTH-1:0] hash_out_6_23;
logic hash_out_valid_filter_6_23;
rule_s_t din_6_23;
rule_s_t din_6_23_r1;
rule_s_t din_6_23_r2;
logic din_valid_6_23;
logic din_valid_6_23_r1;
logic din_valid_6_23_r2;
logic din_ready_6_23;
logic din_almost_full_6_23;
logic [31:0] din_csr_readdata_6_23;
rule_s_t back_data_6_23;
logic    back_valid_6_23;
logic    back_ready_6_23;
logic [RID_WIDTH-1:0] hash_out_6_24;
logic hash_out_valid_filter_6_24;
rule_s_t din_6_24;
rule_s_t din_6_24_r1;
rule_s_t din_6_24_r2;
logic din_valid_6_24;
logic din_valid_6_24_r1;
logic din_valid_6_24_r2;
logic din_ready_6_24;
logic din_almost_full_6_24;
logic [31:0] din_csr_readdata_6_24;
rule_s_t back_data_6_24;
logic    back_valid_6_24;
logic    back_ready_6_24;
logic [RID_WIDTH-1:0] hash_out_6_25;
logic hash_out_valid_filter_6_25;
rule_s_t din_6_25;
rule_s_t din_6_25_r1;
rule_s_t din_6_25_r2;
logic din_valid_6_25;
logic din_valid_6_25_r1;
logic din_valid_6_25_r2;
logic din_ready_6_25;
logic din_almost_full_6_25;
logic [31:0] din_csr_readdata_6_25;
rule_s_t back_data_6_25;
logic    back_valid_6_25;
logic    back_ready_6_25;
logic [RID_WIDTH-1:0] hash_out_6_26;
logic hash_out_valid_filter_6_26;
rule_s_t din_6_26;
rule_s_t din_6_26_r1;
rule_s_t din_6_26_r2;
logic din_valid_6_26;
logic din_valid_6_26_r1;
logic din_valid_6_26_r2;
logic din_ready_6_26;
logic din_almost_full_6_26;
logic [31:0] din_csr_readdata_6_26;
rule_s_t back_data_6_26;
logic    back_valid_6_26;
logic    back_ready_6_26;
logic [RID_WIDTH-1:0] hash_out_6_27;
logic hash_out_valid_filter_6_27;
rule_s_t din_6_27;
rule_s_t din_6_27_r1;
rule_s_t din_6_27_r2;
logic din_valid_6_27;
logic din_valid_6_27_r1;
logic din_valid_6_27_r2;
logic din_ready_6_27;
logic din_almost_full_6_27;
logic [31:0] din_csr_readdata_6_27;
rule_s_t back_data_6_27;
logic    back_valid_6_27;
logic    back_ready_6_27;
logic [RID_WIDTH-1:0] hash_out_6_28;
logic hash_out_valid_filter_6_28;
rule_s_t din_6_28;
rule_s_t din_6_28_r1;
rule_s_t din_6_28_r2;
logic din_valid_6_28;
logic din_valid_6_28_r1;
logic din_valid_6_28_r2;
logic din_ready_6_28;
logic din_almost_full_6_28;
logic [31:0] din_csr_readdata_6_28;
rule_s_t back_data_6_28;
logic    back_valid_6_28;
logic    back_ready_6_28;
logic [RID_WIDTH-1:0] hash_out_6_29;
logic hash_out_valid_filter_6_29;
rule_s_t din_6_29;
rule_s_t din_6_29_r1;
rule_s_t din_6_29_r2;
logic din_valid_6_29;
logic din_valid_6_29_r1;
logic din_valid_6_29_r2;
logic din_ready_6_29;
logic din_almost_full_6_29;
logic [31:0] din_csr_readdata_6_29;
rule_s_t back_data_6_29;
logic    back_valid_6_29;
logic    back_ready_6_29;
logic [RID_WIDTH-1:0] hash_out_6_30;
logic hash_out_valid_filter_6_30;
rule_s_t din_6_30;
rule_s_t din_6_30_r1;
rule_s_t din_6_30_r2;
logic din_valid_6_30;
logic din_valid_6_30_r1;
logic din_valid_6_30_r2;
logic din_ready_6_30;
logic din_almost_full_6_30;
logic [31:0] din_csr_readdata_6_30;
rule_s_t back_data_6_30;
logic    back_valid_6_30;
logic    back_ready_6_30;
logic [RID_WIDTH-1:0] hash_out_6_31;
logic hash_out_valid_filter_6_31;
rule_s_t din_6_31;
rule_s_t din_6_31_r1;
rule_s_t din_6_31_r2;
logic din_valid_6_31;
logic din_valid_6_31_r1;
logic din_valid_6_31_r2;
logic din_ready_6_31;
logic din_almost_full_6_31;
logic [31:0] din_csr_readdata_6_31;
rule_s_t back_data_6_31;
logic    back_valid_6_31;
logic    back_ready_6_31;
logic [RID_WIDTH-1:0] hash_out_7_0;
logic hash_out_valid_filter_7_0;
rule_s_t din_7_0;
rule_s_t din_7_0_r1;
rule_s_t din_7_0_r2;
logic din_valid_7_0;
logic din_valid_7_0_r1;
logic din_valid_7_0_r2;
logic din_ready_7_0;
logic din_almost_full_7_0;
logic [31:0] din_csr_readdata_7_0;
rule_s_t back_data_7_0;
logic    back_valid_7_0;
logic    back_ready_7_0;
logic [RID_WIDTH-1:0] hash_out_7_1;
logic hash_out_valid_filter_7_1;
rule_s_t din_7_1;
rule_s_t din_7_1_r1;
rule_s_t din_7_1_r2;
logic din_valid_7_1;
logic din_valid_7_1_r1;
logic din_valid_7_1_r2;
logic din_ready_7_1;
logic din_almost_full_7_1;
logic [31:0] din_csr_readdata_7_1;
rule_s_t back_data_7_1;
logic    back_valid_7_1;
logic    back_ready_7_1;
logic [RID_WIDTH-1:0] hash_out_7_2;
logic hash_out_valid_filter_7_2;
rule_s_t din_7_2;
rule_s_t din_7_2_r1;
rule_s_t din_7_2_r2;
logic din_valid_7_2;
logic din_valid_7_2_r1;
logic din_valid_7_2_r2;
logic din_ready_7_2;
logic din_almost_full_7_2;
logic [31:0] din_csr_readdata_7_2;
rule_s_t back_data_7_2;
logic    back_valid_7_2;
logic    back_ready_7_2;
logic [RID_WIDTH-1:0] hash_out_7_3;
logic hash_out_valid_filter_7_3;
rule_s_t din_7_3;
rule_s_t din_7_3_r1;
rule_s_t din_7_3_r2;
logic din_valid_7_3;
logic din_valid_7_3_r1;
logic din_valid_7_3_r2;
logic din_ready_7_3;
logic din_almost_full_7_3;
logic [31:0] din_csr_readdata_7_3;
rule_s_t back_data_7_3;
logic    back_valid_7_3;
logic    back_ready_7_3;
logic [RID_WIDTH-1:0] hash_out_7_4;
logic hash_out_valid_filter_7_4;
rule_s_t din_7_4;
rule_s_t din_7_4_r1;
rule_s_t din_7_4_r2;
logic din_valid_7_4;
logic din_valid_7_4_r1;
logic din_valid_7_4_r2;
logic din_ready_7_4;
logic din_almost_full_7_4;
logic [31:0] din_csr_readdata_7_4;
rule_s_t back_data_7_4;
logic    back_valid_7_4;
logic    back_ready_7_4;
logic [RID_WIDTH-1:0] hash_out_7_5;
logic hash_out_valid_filter_7_5;
rule_s_t din_7_5;
rule_s_t din_7_5_r1;
rule_s_t din_7_5_r2;
logic din_valid_7_5;
logic din_valid_7_5_r1;
logic din_valid_7_5_r2;
logic din_ready_7_5;
logic din_almost_full_7_5;
logic [31:0] din_csr_readdata_7_5;
rule_s_t back_data_7_5;
logic    back_valid_7_5;
logic    back_ready_7_5;
logic [RID_WIDTH-1:0] hash_out_7_6;
logic hash_out_valid_filter_7_6;
rule_s_t din_7_6;
rule_s_t din_7_6_r1;
rule_s_t din_7_6_r2;
logic din_valid_7_6;
logic din_valid_7_6_r1;
logic din_valid_7_6_r2;
logic din_ready_7_6;
logic din_almost_full_7_6;
logic [31:0] din_csr_readdata_7_6;
rule_s_t back_data_7_6;
logic    back_valid_7_6;
logic    back_ready_7_6;
logic [RID_WIDTH-1:0] hash_out_7_7;
logic hash_out_valid_filter_7_7;
rule_s_t din_7_7;
rule_s_t din_7_7_r1;
rule_s_t din_7_7_r2;
logic din_valid_7_7;
logic din_valid_7_7_r1;
logic din_valid_7_7_r2;
logic din_ready_7_7;
logic din_almost_full_7_7;
logic [31:0] din_csr_readdata_7_7;
rule_s_t back_data_7_7;
logic    back_valid_7_7;
logic    back_ready_7_7;
logic [RID_WIDTH-1:0] hash_out_7_8;
logic hash_out_valid_filter_7_8;
rule_s_t din_7_8;
rule_s_t din_7_8_r1;
rule_s_t din_7_8_r2;
logic din_valid_7_8;
logic din_valid_7_8_r1;
logic din_valid_7_8_r2;
logic din_ready_7_8;
logic din_almost_full_7_8;
logic [31:0] din_csr_readdata_7_8;
rule_s_t back_data_7_8;
logic    back_valid_7_8;
logic    back_ready_7_8;
logic [RID_WIDTH-1:0] hash_out_7_9;
logic hash_out_valid_filter_7_9;
rule_s_t din_7_9;
rule_s_t din_7_9_r1;
rule_s_t din_7_9_r2;
logic din_valid_7_9;
logic din_valid_7_9_r1;
logic din_valid_7_9_r2;
logic din_ready_7_9;
logic din_almost_full_7_9;
logic [31:0] din_csr_readdata_7_9;
rule_s_t back_data_7_9;
logic    back_valid_7_9;
logic    back_ready_7_9;
logic [RID_WIDTH-1:0] hash_out_7_10;
logic hash_out_valid_filter_7_10;
rule_s_t din_7_10;
rule_s_t din_7_10_r1;
rule_s_t din_7_10_r2;
logic din_valid_7_10;
logic din_valid_7_10_r1;
logic din_valid_7_10_r2;
logic din_ready_7_10;
logic din_almost_full_7_10;
logic [31:0] din_csr_readdata_7_10;
rule_s_t back_data_7_10;
logic    back_valid_7_10;
logic    back_ready_7_10;
logic [RID_WIDTH-1:0] hash_out_7_11;
logic hash_out_valid_filter_7_11;
rule_s_t din_7_11;
rule_s_t din_7_11_r1;
rule_s_t din_7_11_r2;
logic din_valid_7_11;
logic din_valid_7_11_r1;
logic din_valid_7_11_r2;
logic din_ready_7_11;
logic din_almost_full_7_11;
logic [31:0] din_csr_readdata_7_11;
rule_s_t back_data_7_11;
logic    back_valid_7_11;
logic    back_ready_7_11;
logic [RID_WIDTH-1:0] hash_out_7_12;
logic hash_out_valid_filter_7_12;
rule_s_t din_7_12;
rule_s_t din_7_12_r1;
rule_s_t din_7_12_r2;
logic din_valid_7_12;
logic din_valid_7_12_r1;
logic din_valid_7_12_r2;
logic din_ready_7_12;
logic din_almost_full_7_12;
logic [31:0] din_csr_readdata_7_12;
rule_s_t back_data_7_12;
logic    back_valid_7_12;
logic    back_ready_7_12;
logic [RID_WIDTH-1:0] hash_out_7_13;
logic hash_out_valid_filter_7_13;
rule_s_t din_7_13;
rule_s_t din_7_13_r1;
rule_s_t din_7_13_r2;
logic din_valid_7_13;
logic din_valid_7_13_r1;
logic din_valid_7_13_r2;
logic din_ready_7_13;
logic din_almost_full_7_13;
logic [31:0] din_csr_readdata_7_13;
rule_s_t back_data_7_13;
logic    back_valid_7_13;
logic    back_ready_7_13;
logic [RID_WIDTH-1:0] hash_out_7_14;
logic hash_out_valid_filter_7_14;
rule_s_t din_7_14;
rule_s_t din_7_14_r1;
rule_s_t din_7_14_r2;
logic din_valid_7_14;
logic din_valid_7_14_r1;
logic din_valid_7_14_r2;
logic din_ready_7_14;
logic din_almost_full_7_14;
logic [31:0] din_csr_readdata_7_14;
rule_s_t back_data_7_14;
logic    back_valid_7_14;
logic    back_ready_7_14;
logic [RID_WIDTH-1:0] hash_out_7_15;
logic hash_out_valid_filter_7_15;
rule_s_t din_7_15;
rule_s_t din_7_15_r1;
rule_s_t din_7_15_r2;
logic din_valid_7_15;
logic din_valid_7_15_r1;
logic din_valid_7_15_r2;
logic din_ready_7_15;
logic din_almost_full_7_15;
logic [31:0] din_csr_readdata_7_15;
rule_s_t back_data_7_15;
logic    back_valid_7_15;
logic    back_ready_7_15;
logic [RID_WIDTH-1:0] hash_out_7_16;
logic hash_out_valid_filter_7_16;
rule_s_t din_7_16;
rule_s_t din_7_16_r1;
rule_s_t din_7_16_r2;
logic din_valid_7_16;
logic din_valid_7_16_r1;
logic din_valid_7_16_r2;
logic din_ready_7_16;
logic din_almost_full_7_16;
logic [31:0] din_csr_readdata_7_16;
rule_s_t back_data_7_16;
logic    back_valid_7_16;
logic    back_ready_7_16;
logic [RID_WIDTH-1:0] hash_out_7_17;
logic hash_out_valid_filter_7_17;
rule_s_t din_7_17;
rule_s_t din_7_17_r1;
rule_s_t din_7_17_r2;
logic din_valid_7_17;
logic din_valid_7_17_r1;
logic din_valid_7_17_r2;
logic din_ready_7_17;
logic din_almost_full_7_17;
logic [31:0] din_csr_readdata_7_17;
rule_s_t back_data_7_17;
logic    back_valid_7_17;
logic    back_ready_7_17;
logic [RID_WIDTH-1:0] hash_out_7_18;
logic hash_out_valid_filter_7_18;
rule_s_t din_7_18;
rule_s_t din_7_18_r1;
rule_s_t din_7_18_r2;
logic din_valid_7_18;
logic din_valid_7_18_r1;
logic din_valid_7_18_r2;
logic din_ready_7_18;
logic din_almost_full_7_18;
logic [31:0] din_csr_readdata_7_18;
rule_s_t back_data_7_18;
logic    back_valid_7_18;
logic    back_ready_7_18;
logic [RID_WIDTH-1:0] hash_out_7_19;
logic hash_out_valid_filter_7_19;
rule_s_t din_7_19;
rule_s_t din_7_19_r1;
rule_s_t din_7_19_r2;
logic din_valid_7_19;
logic din_valid_7_19_r1;
logic din_valid_7_19_r2;
logic din_ready_7_19;
logic din_almost_full_7_19;
logic [31:0] din_csr_readdata_7_19;
rule_s_t back_data_7_19;
logic    back_valid_7_19;
logic    back_ready_7_19;
logic [RID_WIDTH-1:0] hash_out_7_20;
logic hash_out_valid_filter_7_20;
rule_s_t din_7_20;
rule_s_t din_7_20_r1;
rule_s_t din_7_20_r2;
logic din_valid_7_20;
logic din_valid_7_20_r1;
logic din_valid_7_20_r2;
logic din_ready_7_20;
logic din_almost_full_7_20;
logic [31:0] din_csr_readdata_7_20;
rule_s_t back_data_7_20;
logic    back_valid_7_20;
logic    back_ready_7_20;
logic [RID_WIDTH-1:0] hash_out_7_21;
logic hash_out_valid_filter_7_21;
rule_s_t din_7_21;
rule_s_t din_7_21_r1;
rule_s_t din_7_21_r2;
logic din_valid_7_21;
logic din_valid_7_21_r1;
logic din_valid_7_21_r2;
logic din_ready_7_21;
logic din_almost_full_7_21;
logic [31:0] din_csr_readdata_7_21;
rule_s_t back_data_7_21;
logic    back_valid_7_21;
logic    back_ready_7_21;
logic [RID_WIDTH-1:0] hash_out_7_22;
logic hash_out_valid_filter_7_22;
rule_s_t din_7_22;
rule_s_t din_7_22_r1;
rule_s_t din_7_22_r2;
logic din_valid_7_22;
logic din_valid_7_22_r1;
logic din_valid_7_22_r2;
logic din_ready_7_22;
logic din_almost_full_7_22;
logic [31:0] din_csr_readdata_7_22;
rule_s_t back_data_7_22;
logic    back_valid_7_22;
logic    back_ready_7_22;
logic [RID_WIDTH-1:0] hash_out_7_23;
logic hash_out_valid_filter_7_23;
rule_s_t din_7_23;
rule_s_t din_7_23_r1;
rule_s_t din_7_23_r2;
logic din_valid_7_23;
logic din_valid_7_23_r1;
logic din_valid_7_23_r2;
logic din_ready_7_23;
logic din_almost_full_7_23;
logic [31:0] din_csr_readdata_7_23;
rule_s_t back_data_7_23;
logic    back_valid_7_23;
logic    back_ready_7_23;
logic [RID_WIDTH-1:0] hash_out_7_24;
logic hash_out_valid_filter_7_24;
rule_s_t din_7_24;
rule_s_t din_7_24_r1;
rule_s_t din_7_24_r2;
logic din_valid_7_24;
logic din_valid_7_24_r1;
logic din_valid_7_24_r2;
logic din_ready_7_24;
logic din_almost_full_7_24;
logic [31:0] din_csr_readdata_7_24;
rule_s_t back_data_7_24;
logic    back_valid_7_24;
logic    back_ready_7_24;
logic [RID_WIDTH-1:0] hash_out_7_25;
logic hash_out_valid_filter_7_25;
rule_s_t din_7_25;
rule_s_t din_7_25_r1;
rule_s_t din_7_25_r2;
logic din_valid_7_25;
logic din_valid_7_25_r1;
logic din_valid_7_25_r2;
logic din_ready_7_25;
logic din_almost_full_7_25;
logic [31:0] din_csr_readdata_7_25;
rule_s_t back_data_7_25;
logic    back_valid_7_25;
logic    back_ready_7_25;
logic [RID_WIDTH-1:0] hash_out_7_26;
logic hash_out_valid_filter_7_26;
rule_s_t din_7_26;
rule_s_t din_7_26_r1;
rule_s_t din_7_26_r2;
logic din_valid_7_26;
logic din_valid_7_26_r1;
logic din_valid_7_26_r2;
logic din_ready_7_26;
logic din_almost_full_7_26;
logic [31:0] din_csr_readdata_7_26;
rule_s_t back_data_7_26;
logic    back_valid_7_26;
logic    back_ready_7_26;
logic [RID_WIDTH-1:0] hash_out_7_27;
logic hash_out_valid_filter_7_27;
rule_s_t din_7_27;
rule_s_t din_7_27_r1;
rule_s_t din_7_27_r2;
logic din_valid_7_27;
logic din_valid_7_27_r1;
logic din_valid_7_27_r2;
logic din_ready_7_27;
logic din_almost_full_7_27;
logic [31:0] din_csr_readdata_7_27;
rule_s_t back_data_7_27;
logic    back_valid_7_27;
logic    back_ready_7_27;
logic [RID_WIDTH-1:0] hash_out_7_28;
logic hash_out_valid_filter_7_28;
rule_s_t din_7_28;
rule_s_t din_7_28_r1;
rule_s_t din_7_28_r2;
logic din_valid_7_28;
logic din_valid_7_28_r1;
logic din_valid_7_28_r2;
logic din_ready_7_28;
logic din_almost_full_7_28;
logic [31:0] din_csr_readdata_7_28;
rule_s_t back_data_7_28;
logic    back_valid_7_28;
logic    back_ready_7_28;
logic [RID_WIDTH-1:0] hash_out_7_29;
logic hash_out_valid_filter_7_29;
rule_s_t din_7_29;
rule_s_t din_7_29_r1;
rule_s_t din_7_29_r2;
logic din_valid_7_29;
logic din_valid_7_29_r1;
logic din_valid_7_29_r2;
logic din_ready_7_29;
logic din_almost_full_7_29;
logic [31:0] din_csr_readdata_7_29;
rule_s_t back_data_7_29;
logic    back_valid_7_29;
logic    back_ready_7_29;
logic [RID_WIDTH-1:0] hash_out_7_30;
logic hash_out_valid_filter_7_30;
rule_s_t din_7_30;
rule_s_t din_7_30_r1;
rule_s_t din_7_30_r2;
logic din_valid_7_30;
logic din_valid_7_30_r1;
logic din_valid_7_30_r2;
logic din_ready_7_30;
logic din_almost_full_7_30;
logic [31:0] din_csr_readdata_7_30;
rule_s_t back_data_7_30;
logic    back_valid_7_30;
logic    back_ready_7_30;
logic [RID_WIDTH-1:0] hash_out_7_31;
logic hash_out_valid_filter_7_31;
rule_s_t din_7_31;
rule_s_t din_7_31_r1;
rule_s_t din_7_31_r2;
logic din_valid_7_31;
logic din_valid_7_31_r1;
logic din_valid_7_31_r2;
logic din_ready_7_31;
logic din_almost_full_7_31;
logic [31:0] din_csr_readdata_7_31;
rule_s_t back_data_7_31;
logic    back_valid_7_31;
logic    back_ready_7_31;

logic out_new_pkt;

assign piped_pkt_data_swap[7+0*8:0+0*8] = piped_pkt_data[FP_DWIDTH-1-0*8:FP_DWIDTH-8-0*8];
assign piped_pkt_data_swap[7+1*8:0+1*8] = piped_pkt_data[FP_DWIDTH-1-1*8:FP_DWIDTH-8-1*8];
assign piped_pkt_data_swap[7+2*8:0+2*8] = piped_pkt_data[FP_DWIDTH-1-2*8:FP_DWIDTH-8-2*8];
assign piped_pkt_data_swap[7+3*8:0+3*8] = piped_pkt_data[FP_DWIDTH-1-3*8:FP_DWIDTH-8-3*8];
assign piped_pkt_data_swap[7+4*8:0+4*8] = piped_pkt_data[FP_DWIDTH-1-4*8:FP_DWIDTH-8-4*8];
assign piped_pkt_data_swap[7+5*8:0+5*8] = piped_pkt_data[FP_DWIDTH-1-5*8:FP_DWIDTH-8-5*8];
assign piped_pkt_data_swap[7+6*8:0+6*8] = piped_pkt_data[FP_DWIDTH-1-6*8:FP_DWIDTH-8-6*8];
assign piped_pkt_data_swap[7+7*8:0+7*8] = piped_pkt_data[FP_DWIDTH-1-7*8:FP_DWIDTH-8-7*8];
assign piped_pkt_data_swap[7+8*8:0+8*8] = piped_pkt_data[FP_DWIDTH-1-8*8:FP_DWIDTH-8-8*8];
assign piped_pkt_data_swap[7+9*8:0+9*8] = piped_pkt_data[FP_DWIDTH-1-9*8:FP_DWIDTH-8-9*8];
assign piped_pkt_data_swap[7+10*8:0+10*8] = piped_pkt_data[FP_DWIDTH-1-10*8:FP_DWIDTH-8-10*8];
assign piped_pkt_data_swap[7+11*8:0+11*8] = piped_pkt_data[FP_DWIDTH-1-11*8:FP_DWIDTH-8-11*8];
assign piped_pkt_data_swap[7+12*8:0+12*8] = piped_pkt_data[FP_DWIDTH-1-12*8:FP_DWIDTH-8-12*8];
assign piped_pkt_data_swap[7+13*8:0+13*8] = piped_pkt_data[FP_DWIDTH-1-13*8:FP_DWIDTH-8-13*8];
assign piped_pkt_data_swap[7+14*8:0+14*8] = piped_pkt_data[FP_DWIDTH-1-14*8:FP_DWIDTH-8-14*8];
assign piped_pkt_data_swap[7+15*8:0+15*8] = piped_pkt_data[FP_DWIDTH-1-15*8:FP_DWIDTH-8-15*8];
assign piped_pkt_data_swap[7+16*8:0+16*8] = piped_pkt_data[FP_DWIDTH-1-16*8:FP_DWIDTH-8-16*8];
assign piped_pkt_data_swap[7+17*8:0+17*8] = piped_pkt_data[FP_DWIDTH-1-17*8:FP_DWIDTH-8-17*8];
assign piped_pkt_data_swap[7+18*8:0+18*8] = piped_pkt_data[FP_DWIDTH-1-18*8:FP_DWIDTH-8-18*8];
assign piped_pkt_data_swap[7+19*8:0+19*8] = piped_pkt_data[FP_DWIDTH-1-19*8:FP_DWIDTH-8-19*8];
assign piped_pkt_data_swap[7+20*8:0+20*8] = piped_pkt_data[FP_DWIDTH-1-20*8:FP_DWIDTH-8-20*8];
assign piped_pkt_data_swap[7+21*8:0+21*8] = piped_pkt_data[FP_DWIDTH-1-21*8:FP_DWIDTH-8-21*8];
assign piped_pkt_data_swap[7+22*8:0+22*8] = piped_pkt_data[FP_DWIDTH-1-22*8:FP_DWIDTH-8-22*8];
assign piped_pkt_data_swap[7+23*8:0+23*8] = piped_pkt_data[FP_DWIDTH-1-23*8:FP_DWIDTH-8-23*8];
assign piped_pkt_data_swap[7+24*8:0+24*8] = piped_pkt_data[FP_DWIDTH-1-24*8:FP_DWIDTH-8-24*8];
assign piped_pkt_data_swap[7+25*8:0+25*8] = piped_pkt_data[FP_DWIDTH-1-25*8:FP_DWIDTH-8-25*8];
assign piped_pkt_data_swap[7+26*8:0+26*8] = piped_pkt_data[FP_DWIDTH-1-26*8:FP_DWIDTH-8-26*8];
assign piped_pkt_data_swap[7+27*8:0+27*8] = piped_pkt_data[FP_DWIDTH-1-27*8:FP_DWIDTH-8-27*8];
assign piped_pkt_data_swap[7+28*8:0+28*8] = piped_pkt_data[FP_DWIDTH-1-28*8:FP_DWIDTH-8-28*8];
assign piped_pkt_data_swap[7+29*8:0+29*8] = piped_pkt_data[FP_DWIDTH-1-29*8:FP_DWIDTH-8-29*8];
assign piped_pkt_data_swap[7+30*8:0+30*8] = piped_pkt_data[FP_DWIDTH-1-30*8:FP_DWIDTH-8-30*8];
assign piped_pkt_data_swap[7+31*8:0+31*8] = piped_pkt_data[FP_DWIDTH-1-31*8:FP_DWIDTH-8-31*8];

//Insert retiming register for better timing
always @ (posedge front_clk) begin
    if(front_rst)begin
        piped_pkt_almost_full <= 0;
    end else begin
        piped_pkt_almost_full <=   din_almost_full_0_0 |  din_almost_full_0_1 |  din_almost_full_0_2 |  din_almost_full_0_3 |  din_almost_full_0_4 |  din_almost_full_0_5 |  din_almost_full_0_6 |  din_almost_full_0_7 |  din_almost_full_0_8 |  din_almost_full_0_9 |  din_almost_full_0_10 |  din_almost_full_0_11 |  din_almost_full_0_12 |  din_almost_full_0_13 |  din_almost_full_0_14 |  din_almost_full_0_15 |  din_almost_full_0_16 |  din_almost_full_0_17 |  din_almost_full_0_18 |  din_almost_full_0_19 |  din_almost_full_0_20 |  din_almost_full_0_21 |  din_almost_full_0_22 |  din_almost_full_0_23 |  din_almost_full_0_24 |  din_almost_full_0_25 |  din_almost_full_0_26 |  din_almost_full_0_27 |  din_almost_full_0_28 |  din_almost_full_0_29 |  din_almost_full_0_30 |  din_almost_full_0_31 |    din_almost_full_1_0 |  din_almost_full_1_1 |  din_almost_full_1_2 |  din_almost_full_1_3 |  din_almost_full_1_4 |  din_almost_full_1_5 |  din_almost_full_1_6 |  din_almost_full_1_7 |  din_almost_full_1_8 |  din_almost_full_1_9 |  din_almost_full_1_10 |  din_almost_full_1_11 |  din_almost_full_1_12 |  din_almost_full_1_13 |  din_almost_full_1_14 |  din_almost_full_1_15 |  din_almost_full_1_16 |  din_almost_full_1_17 |  din_almost_full_1_18 |  din_almost_full_1_19 |  din_almost_full_1_20 |  din_almost_full_1_21 |  din_almost_full_1_22 |  din_almost_full_1_23 |  din_almost_full_1_24 |  din_almost_full_1_25 |  din_almost_full_1_26 |  din_almost_full_1_27 |  din_almost_full_1_28 |  din_almost_full_1_29 |  din_almost_full_1_30 |  din_almost_full_1_31 |    din_almost_full_2_0 |  din_almost_full_2_1 |  din_almost_full_2_2 |  din_almost_full_2_3 |  din_almost_full_2_4 |  din_almost_full_2_5 |  din_almost_full_2_6 |  din_almost_full_2_7 |  din_almost_full_2_8 |  din_almost_full_2_9 |  din_almost_full_2_10 |  din_almost_full_2_11 |  din_almost_full_2_12 |  din_almost_full_2_13 |  din_almost_full_2_14 |  din_almost_full_2_15 |  din_almost_full_2_16 |  din_almost_full_2_17 |  din_almost_full_2_18 |  din_almost_full_2_19 |  din_almost_full_2_20 |  din_almost_full_2_21 |  din_almost_full_2_22 |  din_almost_full_2_23 |  din_almost_full_2_24 |  din_almost_full_2_25 |  din_almost_full_2_26 |  din_almost_full_2_27 |  din_almost_full_2_28 |  din_almost_full_2_29 |  din_almost_full_2_30 |  din_almost_full_2_31 |    din_almost_full_3_0 |  din_almost_full_3_1 |  din_almost_full_3_2 |  din_almost_full_3_3 |  din_almost_full_3_4 |  din_almost_full_3_5 |  din_almost_full_3_6 |  din_almost_full_3_7 |  din_almost_full_3_8 |  din_almost_full_3_9 |  din_almost_full_3_10 |  din_almost_full_3_11 |  din_almost_full_3_12 |  din_almost_full_3_13 |  din_almost_full_3_14 |  din_almost_full_3_15 |  din_almost_full_3_16 |  din_almost_full_3_17 |  din_almost_full_3_18 |  din_almost_full_3_19 |  din_almost_full_3_20 |  din_almost_full_3_21 |  din_almost_full_3_22 |  din_almost_full_3_23 |  din_almost_full_3_24 |  din_almost_full_3_25 |  din_almost_full_3_26 |  din_almost_full_3_27 |  din_almost_full_3_28 |  din_almost_full_3_29 |  din_almost_full_3_30 |  din_almost_full_3_31 |    din_almost_full_4_0 |  din_almost_full_4_1 |  din_almost_full_4_2 |  din_almost_full_4_3 |  din_almost_full_4_4 |  din_almost_full_4_5 |  din_almost_full_4_6 |  din_almost_full_4_7 |  din_almost_full_4_8 |  din_almost_full_4_9 |  din_almost_full_4_10 |  din_almost_full_4_11 |  din_almost_full_4_12 |  din_almost_full_4_13 |  din_almost_full_4_14 |  din_almost_full_4_15 |  din_almost_full_4_16 |  din_almost_full_4_17 |  din_almost_full_4_18 |  din_almost_full_4_19 |  din_almost_full_4_20 |  din_almost_full_4_21 |  din_almost_full_4_22 |  din_almost_full_4_23 |  din_almost_full_4_24 |  din_almost_full_4_25 |  din_almost_full_4_26 |  din_almost_full_4_27 |  din_almost_full_4_28 |  din_almost_full_4_29 |  din_almost_full_4_30 |  din_almost_full_4_31 |    din_almost_full_5_0 |  din_almost_full_5_1 |  din_almost_full_5_2 |  din_almost_full_5_3 |  din_almost_full_5_4 |  din_almost_full_5_5 |  din_almost_full_5_6 |  din_almost_full_5_7 |  din_almost_full_5_8 |  din_almost_full_5_9 |  din_almost_full_5_10 |  din_almost_full_5_11 |  din_almost_full_5_12 |  din_almost_full_5_13 |  din_almost_full_5_14 |  din_almost_full_5_15 |  din_almost_full_5_16 |  din_almost_full_5_17 |  din_almost_full_5_18 |  din_almost_full_5_19 |  din_almost_full_5_20 |  din_almost_full_5_21 |  din_almost_full_5_22 |  din_almost_full_5_23 |  din_almost_full_5_24 |  din_almost_full_5_25 |  din_almost_full_5_26 |  din_almost_full_5_27 |  din_almost_full_5_28 |  din_almost_full_5_29 |  din_almost_full_5_30 |  din_almost_full_5_31 |    din_almost_full_6_0 |  din_almost_full_6_1 |  din_almost_full_6_2 |  din_almost_full_6_3 |  din_almost_full_6_4 |  din_almost_full_6_5 |  din_almost_full_6_6 |  din_almost_full_6_7 |  din_almost_full_6_8 |  din_almost_full_6_9 |  din_almost_full_6_10 |  din_almost_full_6_11 |  din_almost_full_6_12 |  din_almost_full_6_13 |  din_almost_full_6_14 |  din_almost_full_6_15 |  din_almost_full_6_16 |  din_almost_full_6_17 |  din_almost_full_6_18 |  din_almost_full_6_19 |  din_almost_full_6_20 |  din_almost_full_6_21 |  din_almost_full_6_22 |  din_almost_full_6_23 |  din_almost_full_6_24 |  din_almost_full_6_25 |  din_almost_full_6_26 |  din_almost_full_6_27 |  din_almost_full_6_28 |  din_almost_full_6_29 |  din_almost_full_6_30 |  din_almost_full_6_31 |    din_almost_full_7_0 |  din_almost_full_7_1 |  din_almost_full_7_2 |  din_almost_full_7_3 |  din_almost_full_7_4 |  din_almost_full_7_5 |  din_almost_full_7_6 |  din_almost_full_7_7 |  din_almost_full_7_8 |  din_almost_full_7_9 |  din_almost_full_7_10 |  din_almost_full_7_11 |  din_almost_full_7_12 |  din_almost_full_7_13 |  din_almost_full_7_14 |  din_almost_full_7_15 |  din_almost_full_7_16 |  din_almost_full_7_17 |  din_almost_full_7_18 |  din_almost_full_7_19 |  din_almost_full_7_20 |  din_almost_full_7_21 |  din_almost_full_7_22 |  din_almost_full_7_23 |  din_almost_full_7_24 |  din_almost_full_7_25 |  din_almost_full_7_26 |  din_almost_full_7_27 |  din_almost_full_7_28 |  din_almost_full_7_29 |  din_almost_full_7_30 |  din_almost_full_7_31 |   0;
    end
end

//Debug
//always @ (posedge front_clk) begin
//    
//    
//   if (din_almost_full_0_0) begin
//       $display("din_almost_full_0_0");
//   end  
//   if (din_valid_0_0_r2 & !din_ready_0_0)begin
//       $display("overflow din_0_0");
//       $finish;
//   end
//    
//   if (din_almost_full_0_1) begin
//       $display("din_almost_full_0_1");
//   end  
//   if (din_valid_0_1_r2 & !din_ready_0_1)begin
//       $display("overflow din_0_1");
//       $finish;
//   end
//    
//   if (din_almost_full_0_2) begin
//       $display("din_almost_full_0_2");
//   end  
//   if (din_valid_0_2_r2 & !din_ready_0_2)begin
//       $display("overflow din_0_2");
//       $finish;
//   end
//    
//   if (din_almost_full_0_3) begin
//       $display("din_almost_full_0_3");
//   end  
//   if (din_valid_0_3_r2 & !din_ready_0_3)begin
//       $display("overflow din_0_3");
//       $finish;
//   end
//    
//   if (din_almost_full_0_4) begin
//       $display("din_almost_full_0_4");
//   end  
//   if (din_valid_0_4_r2 & !din_ready_0_4)begin
//       $display("overflow din_0_4");
//       $finish;
//   end
//    
//   if (din_almost_full_0_5) begin
//       $display("din_almost_full_0_5");
//   end  
//   if (din_valid_0_5_r2 & !din_ready_0_5)begin
//       $display("overflow din_0_5");
//       $finish;
//   end
//    
//   if (din_almost_full_0_6) begin
//       $display("din_almost_full_0_6");
//   end  
//   if (din_valid_0_6_r2 & !din_ready_0_6)begin
//       $display("overflow din_0_6");
//       $finish;
//   end
//    
//   if (din_almost_full_0_7) begin
//       $display("din_almost_full_0_7");
//   end  
//   if (din_valid_0_7_r2 & !din_ready_0_7)begin
//       $display("overflow din_0_7");
//       $finish;
//   end
//    
//   if (din_almost_full_0_8) begin
//       $display("din_almost_full_0_8");
//   end  
//   if (din_valid_0_8_r2 & !din_ready_0_8)begin
//       $display("overflow din_0_8");
//       $finish;
//   end
//    
//   if (din_almost_full_0_9) begin
//       $display("din_almost_full_0_9");
//   end  
//   if (din_valid_0_9_r2 & !din_ready_0_9)begin
//       $display("overflow din_0_9");
//       $finish;
//   end
//    
//   if (din_almost_full_0_10) begin
//       $display("din_almost_full_0_10");
//   end  
//   if (din_valid_0_10_r2 & !din_ready_0_10)begin
//       $display("overflow din_0_10");
//       $finish;
//   end
//    
//   if (din_almost_full_0_11) begin
//       $display("din_almost_full_0_11");
//   end  
//   if (din_valid_0_11_r2 & !din_ready_0_11)begin
//       $display("overflow din_0_11");
//       $finish;
//   end
//    
//   if (din_almost_full_0_12) begin
//       $display("din_almost_full_0_12");
//   end  
//   if (din_valid_0_12_r2 & !din_ready_0_12)begin
//       $display("overflow din_0_12");
//       $finish;
//   end
//    
//   if (din_almost_full_0_13) begin
//       $display("din_almost_full_0_13");
//   end  
//   if (din_valid_0_13_r2 & !din_ready_0_13)begin
//       $display("overflow din_0_13");
//       $finish;
//   end
//    
//   if (din_almost_full_0_14) begin
//       $display("din_almost_full_0_14");
//   end  
//   if (din_valid_0_14_r2 & !din_ready_0_14)begin
//       $display("overflow din_0_14");
//       $finish;
//   end
//    
//   if (din_almost_full_0_15) begin
//       $display("din_almost_full_0_15");
//   end  
//   if (din_valid_0_15_r2 & !din_ready_0_15)begin
//       $display("overflow din_0_15");
//       $finish;
//   end
//    
//   if (din_almost_full_0_16) begin
//       $display("din_almost_full_0_16");
//   end  
//   if (din_valid_0_16_r2 & !din_ready_0_16)begin
//       $display("overflow din_0_16");
//       $finish;
//   end
//    
//   if (din_almost_full_0_17) begin
//       $display("din_almost_full_0_17");
//   end  
//   if (din_valid_0_17_r2 & !din_ready_0_17)begin
//       $display("overflow din_0_17");
//       $finish;
//   end
//    
//   if (din_almost_full_0_18) begin
//       $display("din_almost_full_0_18");
//   end  
//   if (din_valid_0_18_r2 & !din_ready_0_18)begin
//       $display("overflow din_0_18");
//       $finish;
//   end
//    
//   if (din_almost_full_0_19) begin
//       $display("din_almost_full_0_19");
//   end  
//   if (din_valid_0_19_r2 & !din_ready_0_19)begin
//       $display("overflow din_0_19");
//       $finish;
//   end
//    
//   if (din_almost_full_0_20) begin
//       $display("din_almost_full_0_20");
//   end  
//   if (din_valid_0_20_r2 & !din_ready_0_20)begin
//       $display("overflow din_0_20");
//       $finish;
//   end
//    
//   if (din_almost_full_0_21) begin
//       $display("din_almost_full_0_21");
//   end  
//   if (din_valid_0_21_r2 & !din_ready_0_21)begin
//       $display("overflow din_0_21");
//       $finish;
//   end
//    
//   if (din_almost_full_0_22) begin
//       $display("din_almost_full_0_22");
//   end  
//   if (din_valid_0_22_r2 & !din_ready_0_22)begin
//       $display("overflow din_0_22");
//       $finish;
//   end
//    
//   if (din_almost_full_0_23) begin
//       $display("din_almost_full_0_23");
//   end  
//   if (din_valid_0_23_r2 & !din_ready_0_23)begin
//       $display("overflow din_0_23");
//       $finish;
//   end
//    
//   if (din_almost_full_0_24) begin
//       $display("din_almost_full_0_24");
//   end  
//   if (din_valid_0_24_r2 & !din_ready_0_24)begin
//       $display("overflow din_0_24");
//       $finish;
//   end
//    
//   if (din_almost_full_0_25) begin
//       $display("din_almost_full_0_25");
//   end  
//   if (din_valid_0_25_r2 & !din_ready_0_25)begin
//       $display("overflow din_0_25");
//       $finish;
//   end
//    
//   if (din_almost_full_0_26) begin
//       $display("din_almost_full_0_26");
//   end  
//   if (din_valid_0_26_r2 & !din_ready_0_26)begin
//       $display("overflow din_0_26");
//       $finish;
//   end
//    
//   if (din_almost_full_0_27) begin
//       $display("din_almost_full_0_27");
//   end  
//   if (din_valid_0_27_r2 & !din_ready_0_27)begin
//       $display("overflow din_0_27");
//       $finish;
//   end
//    
//   if (din_almost_full_0_28) begin
//       $display("din_almost_full_0_28");
//   end  
//   if (din_valid_0_28_r2 & !din_ready_0_28)begin
//       $display("overflow din_0_28");
//       $finish;
//   end
//    
//   if (din_almost_full_0_29) begin
//       $display("din_almost_full_0_29");
//   end  
//   if (din_valid_0_29_r2 & !din_ready_0_29)begin
//       $display("overflow din_0_29");
//       $finish;
//   end
//    
//   if (din_almost_full_0_30) begin
//       $display("din_almost_full_0_30");
//   end  
//   if (din_valid_0_30_r2 & !din_ready_0_30)begin
//       $display("overflow din_0_30");
//       $finish;
//   end
//    
//   if (din_almost_full_0_31) begin
//       $display("din_almost_full_0_31");
//   end  
//   if (din_valid_0_31_r2 & !din_ready_0_31)begin
//       $display("overflow din_0_31");
//       $finish;
//   end
//    
//    
//    
//   if (din_almost_full_1_0) begin
//       $display("din_almost_full_1_0");
//   end  
//   if (din_valid_1_0_r2 & !din_ready_1_0)begin
//       $display("overflow din_1_0");
//       $finish;
//   end
//    
//   if (din_almost_full_1_1) begin
//       $display("din_almost_full_1_1");
//   end  
//   if (din_valid_1_1_r2 & !din_ready_1_1)begin
//       $display("overflow din_1_1");
//       $finish;
//   end
//    
//   if (din_almost_full_1_2) begin
//       $display("din_almost_full_1_2");
//   end  
//   if (din_valid_1_2_r2 & !din_ready_1_2)begin
//       $display("overflow din_1_2");
//       $finish;
//   end
//    
//   if (din_almost_full_1_3) begin
//       $display("din_almost_full_1_3");
//   end  
//   if (din_valid_1_3_r2 & !din_ready_1_3)begin
//       $display("overflow din_1_3");
//       $finish;
//   end
//    
//   if (din_almost_full_1_4) begin
//       $display("din_almost_full_1_4");
//   end  
//   if (din_valid_1_4_r2 & !din_ready_1_4)begin
//       $display("overflow din_1_4");
//       $finish;
//   end
//    
//   if (din_almost_full_1_5) begin
//       $display("din_almost_full_1_5");
//   end  
//   if (din_valid_1_5_r2 & !din_ready_1_5)begin
//       $display("overflow din_1_5");
//       $finish;
//   end
//    
//   if (din_almost_full_1_6) begin
//       $display("din_almost_full_1_6");
//   end  
//   if (din_valid_1_6_r2 & !din_ready_1_6)begin
//       $display("overflow din_1_6");
//       $finish;
//   end
//    
//   if (din_almost_full_1_7) begin
//       $display("din_almost_full_1_7");
//   end  
//   if (din_valid_1_7_r2 & !din_ready_1_7)begin
//       $display("overflow din_1_7");
//       $finish;
//   end
//    
//   if (din_almost_full_1_8) begin
//       $display("din_almost_full_1_8");
//   end  
//   if (din_valid_1_8_r2 & !din_ready_1_8)begin
//       $display("overflow din_1_8");
//       $finish;
//   end
//    
//   if (din_almost_full_1_9) begin
//       $display("din_almost_full_1_9");
//   end  
//   if (din_valid_1_9_r2 & !din_ready_1_9)begin
//       $display("overflow din_1_9");
//       $finish;
//   end
//    
//   if (din_almost_full_1_10) begin
//       $display("din_almost_full_1_10");
//   end  
//   if (din_valid_1_10_r2 & !din_ready_1_10)begin
//       $display("overflow din_1_10");
//       $finish;
//   end
//    
//   if (din_almost_full_1_11) begin
//       $display("din_almost_full_1_11");
//   end  
//   if (din_valid_1_11_r2 & !din_ready_1_11)begin
//       $display("overflow din_1_11");
//       $finish;
//   end
//    
//   if (din_almost_full_1_12) begin
//       $display("din_almost_full_1_12");
//   end  
//   if (din_valid_1_12_r2 & !din_ready_1_12)begin
//       $display("overflow din_1_12");
//       $finish;
//   end
//    
//   if (din_almost_full_1_13) begin
//       $display("din_almost_full_1_13");
//   end  
//   if (din_valid_1_13_r2 & !din_ready_1_13)begin
//       $display("overflow din_1_13");
//       $finish;
//   end
//    
//   if (din_almost_full_1_14) begin
//       $display("din_almost_full_1_14");
//   end  
//   if (din_valid_1_14_r2 & !din_ready_1_14)begin
//       $display("overflow din_1_14");
//       $finish;
//   end
//    
//   if (din_almost_full_1_15) begin
//       $display("din_almost_full_1_15");
//   end  
//   if (din_valid_1_15_r2 & !din_ready_1_15)begin
//       $display("overflow din_1_15");
//       $finish;
//   end
//    
//   if (din_almost_full_1_16) begin
//       $display("din_almost_full_1_16");
//   end  
//   if (din_valid_1_16_r2 & !din_ready_1_16)begin
//       $display("overflow din_1_16");
//       $finish;
//   end
//    
//   if (din_almost_full_1_17) begin
//       $display("din_almost_full_1_17");
//   end  
//   if (din_valid_1_17_r2 & !din_ready_1_17)begin
//       $display("overflow din_1_17");
//       $finish;
//   end
//    
//   if (din_almost_full_1_18) begin
//       $display("din_almost_full_1_18");
//   end  
//   if (din_valid_1_18_r2 & !din_ready_1_18)begin
//       $display("overflow din_1_18");
//       $finish;
//   end
//    
//   if (din_almost_full_1_19) begin
//       $display("din_almost_full_1_19");
//   end  
//   if (din_valid_1_19_r2 & !din_ready_1_19)begin
//       $display("overflow din_1_19");
//       $finish;
//   end
//    
//   if (din_almost_full_1_20) begin
//       $display("din_almost_full_1_20");
//   end  
//   if (din_valid_1_20_r2 & !din_ready_1_20)begin
//       $display("overflow din_1_20");
//       $finish;
//   end
//    
//   if (din_almost_full_1_21) begin
//       $display("din_almost_full_1_21");
//   end  
//   if (din_valid_1_21_r2 & !din_ready_1_21)begin
//       $display("overflow din_1_21");
//       $finish;
//   end
//    
//   if (din_almost_full_1_22) begin
//       $display("din_almost_full_1_22");
//   end  
//   if (din_valid_1_22_r2 & !din_ready_1_22)begin
//       $display("overflow din_1_22");
//       $finish;
//   end
//    
//   if (din_almost_full_1_23) begin
//       $display("din_almost_full_1_23");
//   end  
//   if (din_valid_1_23_r2 & !din_ready_1_23)begin
//       $display("overflow din_1_23");
//       $finish;
//   end
//    
//   if (din_almost_full_1_24) begin
//       $display("din_almost_full_1_24");
//   end  
//   if (din_valid_1_24_r2 & !din_ready_1_24)begin
//       $display("overflow din_1_24");
//       $finish;
//   end
//    
//   if (din_almost_full_1_25) begin
//       $display("din_almost_full_1_25");
//   end  
//   if (din_valid_1_25_r2 & !din_ready_1_25)begin
//       $display("overflow din_1_25");
//       $finish;
//   end
//    
//   if (din_almost_full_1_26) begin
//       $display("din_almost_full_1_26");
//   end  
//   if (din_valid_1_26_r2 & !din_ready_1_26)begin
//       $display("overflow din_1_26");
//       $finish;
//   end
//    
//   if (din_almost_full_1_27) begin
//       $display("din_almost_full_1_27");
//   end  
//   if (din_valid_1_27_r2 & !din_ready_1_27)begin
//       $display("overflow din_1_27");
//       $finish;
//   end
//    
//   if (din_almost_full_1_28) begin
//       $display("din_almost_full_1_28");
//   end  
//   if (din_valid_1_28_r2 & !din_ready_1_28)begin
//       $display("overflow din_1_28");
//       $finish;
//   end
//    
//   if (din_almost_full_1_29) begin
//       $display("din_almost_full_1_29");
//   end  
//   if (din_valid_1_29_r2 & !din_ready_1_29)begin
//       $display("overflow din_1_29");
//       $finish;
//   end
//    
//   if (din_almost_full_1_30) begin
//       $display("din_almost_full_1_30");
//   end  
//   if (din_valid_1_30_r2 & !din_ready_1_30)begin
//       $display("overflow din_1_30");
//       $finish;
//   end
//    
//   if (din_almost_full_1_31) begin
//       $display("din_almost_full_1_31");
//   end  
//   if (din_valid_1_31_r2 & !din_ready_1_31)begin
//       $display("overflow din_1_31");
//       $finish;
//   end
//    
//    
//    
//   if (din_almost_full_2_0) begin
//       $display("din_almost_full_2_0");
//   end  
//   if (din_valid_2_0_r2 & !din_ready_2_0)begin
//       $display("overflow din_2_0");
//       $finish;
//   end
//    
//   if (din_almost_full_2_1) begin
//       $display("din_almost_full_2_1");
//   end  
//   if (din_valid_2_1_r2 & !din_ready_2_1)begin
//       $display("overflow din_2_1");
//       $finish;
//   end
//    
//   if (din_almost_full_2_2) begin
//       $display("din_almost_full_2_2");
//   end  
//   if (din_valid_2_2_r2 & !din_ready_2_2)begin
//       $display("overflow din_2_2");
//       $finish;
//   end
//    
//   if (din_almost_full_2_3) begin
//       $display("din_almost_full_2_3");
//   end  
//   if (din_valid_2_3_r2 & !din_ready_2_3)begin
//       $display("overflow din_2_3");
//       $finish;
//   end
//    
//   if (din_almost_full_2_4) begin
//       $display("din_almost_full_2_4");
//   end  
//   if (din_valid_2_4_r2 & !din_ready_2_4)begin
//       $display("overflow din_2_4");
//       $finish;
//   end
//    
//   if (din_almost_full_2_5) begin
//       $display("din_almost_full_2_5");
//   end  
//   if (din_valid_2_5_r2 & !din_ready_2_5)begin
//       $display("overflow din_2_5");
//       $finish;
//   end
//    
//   if (din_almost_full_2_6) begin
//       $display("din_almost_full_2_6");
//   end  
//   if (din_valid_2_6_r2 & !din_ready_2_6)begin
//       $display("overflow din_2_6");
//       $finish;
//   end
//    
//   if (din_almost_full_2_7) begin
//       $display("din_almost_full_2_7");
//   end  
//   if (din_valid_2_7_r2 & !din_ready_2_7)begin
//       $display("overflow din_2_7");
//       $finish;
//   end
//    
//   if (din_almost_full_2_8) begin
//       $display("din_almost_full_2_8");
//   end  
//   if (din_valid_2_8_r2 & !din_ready_2_8)begin
//       $display("overflow din_2_8");
//       $finish;
//   end
//    
//   if (din_almost_full_2_9) begin
//       $display("din_almost_full_2_9");
//   end  
//   if (din_valid_2_9_r2 & !din_ready_2_9)begin
//       $display("overflow din_2_9");
//       $finish;
//   end
//    
//   if (din_almost_full_2_10) begin
//       $display("din_almost_full_2_10");
//   end  
//   if (din_valid_2_10_r2 & !din_ready_2_10)begin
//       $display("overflow din_2_10");
//       $finish;
//   end
//    
//   if (din_almost_full_2_11) begin
//       $display("din_almost_full_2_11");
//   end  
//   if (din_valid_2_11_r2 & !din_ready_2_11)begin
//       $display("overflow din_2_11");
//       $finish;
//   end
//    
//   if (din_almost_full_2_12) begin
//       $display("din_almost_full_2_12");
//   end  
//   if (din_valid_2_12_r2 & !din_ready_2_12)begin
//       $display("overflow din_2_12");
//       $finish;
//   end
//    
//   if (din_almost_full_2_13) begin
//       $display("din_almost_full_2_13");
//   end  
//   if (din_valid_2_13_r2 & !din_ready_2_13)begin
//       $display("overflow din_2_13");
//       $finish;
//   end
//    
//   if (din_almost_full_2_14) begin
//       $display("din_almost_full_2_14");
//   end  
//   if (din_valid_2_14_r2 & !din_ready_2_14)begin
//       $display("overflow din_2_14");
//       $finish;
//   end
//    
//   if (din_almost_full_2_15) begin
//       $display("din_almost_full_2_15");
//   end  
//   if (din_valid_2_15_r2 & !din_ready_2_15)begin
//       $display("overflow din_2_15");
//       $finish;
//   end
//    
//   if (din_almost_full_2_16) begin
//       $display("din_almost_full_2_16");
//   end  
//   if (din_valid_2_16_r2 & !din_ready_2_16)begin
//       $display("overflow din_2_16");
//       $finish;
//   end
//    
//   if (din_almost_full_2_17) begin
//       $display("din_almost_full_2_17");
//   end  
//   if (din_valid_2_17_r2 & !din_ready_2_17)begin
//       $display("overflow din_2_17");
//       $finish;
//   end
//    
//   if (din_almost_full_2_18) begin
//       $display("din_almost_full_2_18");
//   end  
//   if (din_valid_2_18_r2 & !din_ready_2_18)begin
//       $display("overflow din_2_18");
//       $finish;
//   end
//    
//   if (din_almost_full_2_19) begin
//       $display("din_almost_full_2_19");
//   end  
//   if (din_valid_2_19_r2 & !din_ready_2_19)begin
//       $display("overflow din_2_19");
//       $finish;
//   end
//    
//   if (din_almost_full_2_20) begin
//       $display("din_almost_full_2_20");
//   end  
//   if (din_valid_2_20_r2 & !din_ready_2_20)begin
//       $display("overflow din_2_20");
//       $finish;
//   end
//    
//   if (din_almost_full_2_21) begin
//       $display("din_almost_full_2_21");
//   end  
//   if (din_valid_2_21_r2 & !din_ready_2_21)begin
//       $display("overflow din_2_21");
//       $finish;
//   end
//    
//   if (din_almost_full_2_22) begin
//       $display("din_almost_full_2_22");
//   end  
//   if (din_valid_2_22_r2 & !din_ready_2_22)begin
//       $display("overflow din_2_22");
//       $finish;
//   end
//    
//   if (din_almost_full_2_23) begin
//       $display("din_almost_full_2_23");
//   end  
//   if (din_valid_2_23_r2 & !din_ready_2_23)begin
//       $display("overflow din_2_23");
//       $finish;
//   end
//    
//   if (din_almost_full_2_24) begin
//       $display("din_almost_full_2_24");
//   end  
//   if (din_valid_2_24_r2 & !din_ready_2_24)begin
//       $display("overflow din_2_24");
//       $finish;
//   end
//    
//   if (din_almost_full_2_25) begin
//       $display("din_almost_full_2_25");
//   end  
//   if (din_valid_2_25_r2 & !din_ready_2_25)begin
//       $display("overflow din_2_25");
//       $finish;
//   end
//    
//   if (din_almost_full_2_26) begin
//       $display("din_almost_full_2_26");
//   end  
//   if (din_valid_2_26_r2 & !din_ready_2_26)begin
//       $display("overflow din_2_26");
//       $finish;
//   end
//    
//   if (din_almost_full_2_27) begin
//       $display("din_almost_full_2_27");
//   end  
//   if (din_valid_2_27_r2 & !din_ready_2_27)begin
//       $display("overflow din_2_27");
//       $finish;
//   end
//    
//   if (din_almost_full_2_28) begin
//       $display("din_almost_full_2_28");
//   end  
//   if (din_valid_2_28_r2 & !din_ready_2_28)begin
//       $display("overflow din_2_28");
//       $finish;
//   end
//    
//   if (din_almost_full_2_29) begin
//       $display("din_almost_full_2_29");
//   end  
//   if (din_valid_2_29_r2 & !din_ready_2_29)begin
//       $display("overflow din_2_29");
//       $finish;
//   end
//    
//   if (din_almost_full_2_30) begin
//       $display("din_almost_full_2_30");
//   end  
//   if (din_valid_2_30_r2 & !din_ready_2_30)begin
//       $display("overflow din_2_30");
//       $finish;
//   end
//    
//   if (din_almost_full_2_31) begin
//       $display("din_almost_full_2_31");
//   end  
//   if (din_valid_2_31_r2 & !din_ready_2_31)begin
//       $display("overflow din_2_31");
//       $finish;
//   end
//    
//    
//    
//   if (din_almost_full_3_0) begin
//       $display("din_almost_full_3_0");
//   end  
//   if (din_valid_3_0_r2 & !din_ready_3_0)begin
//       $display("overflow din_3_0");
//       $finish;
//   end
//    
//   if (din_almost_full_3_1) begin
//       $display("din_almost_full_3_1");
//   end  
//   if (din_valid_3_1_r2 & !din_ready_3_1)begin
//       $display("overflow din_3_1");
//       $finish;
//   end
//    
//   if (din_almost_full_3_2) begin
//       $display("din_almost_full_3_2");
//   end  
//   if (din_valid_3_2_r2 & !din_ready_3_2)begin
//       $display("overflow din_3_2");
//       $finish;
//   end
//    
//   if (din_almost_full_3_3) begin
//       $display("din_almost_full_3_3");
//   end  
//   if (din_valid_3_3_r2 & !din_ready_3_3)begin
//       $display("overflow din_3_3");
//       $finish;
//   end
//    
//   if (din_almost_full_3_4) begin
//       $display("din_almost_full_3_4");
//   end  
//   if (din_valid_3_4_r2 & !din_ready_3_4)begin
//       $display("overflow din_3_4");
//       $finish;
//   end
//    
//   if (din_almost_full_3_5) begin
//       $display("din_almost_full_3_5");
//   end  
//   if (din_valid_3_5_r2 & !din_ready_3_5)begin
//       $display("overflow din_3_5");
//       $finish;
//   end
//    
//   if (din_almost_full_3_6) begin
//       $display("din_almost_full_3_6");
//   end  
//   if (din_valid_3_6_r2 & !din_ready_3_6)begin
//       $display("overflow din_3_6");
//       $finish;
//   end
//    
//   if (din_almost_full_3_7) begin
//       $display("din_almost_full_3_7");
//   end  
//   if (din_valid_3_7_r2 & !din_ready_3_7)begin
//       $display("overflow din_3_7");
//       $finish;
//   end
//    
//   if (din_almost_full_3_8) begin
//       $display("din_almost_full_3_8");
//   end  
//   if (din_valid_3_8_r2 & !din_ready_3_8)begin
//       $display("overflow din_3_8");
//       $finish;
//   end
//    
//   if (din_almost_full_3_9) begin
//       $display("din_almost_full_3_9");
//   end  
//   if (din_valid_3_9_r2 & !din_ready_3_9)begin
//       $display("overflow din_3_9");
//       $finish;
//   end
//    
//   if (din_almost_full_3_10) begin
//       $display("din_almost_full_3_10");
//   end  
//   if (din_valid_3_10_r2 & !din_ready_3_10)begin
//       $display("overflow din_3_10");
//       $finish;
//   end
//    
//   if (din_almost_full_3_11) begin
//       $display("din_almost_full_3_11");
//   end  
//   if (din_valid_3_11_r2 & !din_ready_3_11)begin
//       $display("overflow din_3_11");
//       $finish;
//   end
//    
//   if (din_almost_full_3_12) begin
//       $display("din_almost_full_3_12");
//   end  
//   if (din_valid_3_12_r2 & !din_ready_3_12)begin
//       $display("overflow din_3_12");
//       $finish;
//   end
//    
//   if (din_almost_full_3_13) begin
//       $display("din_almost_full_3_13");
//   end  
//   if (din_valid_3_13_r2 & !din_ready_3_13)begin
//       $display("overflow din_3_13");
//       $finish;
//   end
//    
//   if (din_almost_full_3_14) begin
//       $display("din_almost_full_3_14");
//   end  
//   if (din_valid_3_14_r2 & !din_ready_3_14)begin
//       $display("overflow din_3_14");
//       $finish;
//   end
//    
//   if (din_almost_full_3_15) begin
//       $display("din_almost_full_3_15");
//   end  
//   if (din_valid_3_15_r2 & !din_ready_3_15)begin
//       $display("overflow din_3_15");
//       $finish;
//   end
//    
//   if (din_almost_full_3_16) begin
//       $display("din_almost_full_3_16");
//   end  
//   if (din_valid_3_16_r2 & !din_ready_3_16)begin
//       $display("overflow din_3_16");
//       $finish;
//   end
//    
//   if (din_almost_full_3_17) begin
//       $display("din_almost_full_3_17");
//   end  
//   if (din_valid_3_17_r2 & !din_ready_3_17)begin
//       $display("overflow din_3_17");
//       $finish;
//   end
//    
//   if (din_almost_full_3_18) begin
//       $display("din_almost_full_3_18");
//   end  
//   if (din_valid_3_18_r2 & !din_ready_3_18)begin
//       $display("overflow din_3_18");
//       $finish;
//   end
//    
//   if (din_almost_full_3_19) begin
//       $display("din_almost_full_3_19");
//   end  
//   if (din_valid_3_19_r2 & !din_ready_3_19)begin
//       $display("overflow din_3_19");
//       $finish;
//   end
//    
//   if (din_almost_full_3_20) begin
//       $display("din_almost_full_3_20");
//   end  
//   if (din_valid_3_20_r2 & !din_ready_3_20)begin
//       $display("overflow din_3_20");
//       $finish;
//   end
//    
//   if (din_almost_full_3_21) begin
//       $display("din_almost_full_3_21");
//   end  
//   if (din_valid_3_21_r2 & !din_ready_3_21)begin
//       $display("overflow din_3_21");
//       $finish;
//   end
//    
//   if (din_almost_full_3_22) begin
//       $display("din_almost_full_3_22");
//   end  
//   if (din_valid_3_22_r2 & !din_ready_3_22)begin
//       $display("overflow din_3_22");
//       $finish;
//   end
//    
//   if (din_almost_full_3_23) begin
//       $display("din_almost_full_3_23");
//   end  
//   if (din_valid_3_23_r2 & !din_ready_3_23)begin
//       $display("overflow din_3_23");
//       $finish;
//   end
//    
//   if (din_almost_full_3_24) begin
//       $display("din_almost_full_3_24");
//   end  
//   if (din_valid_3_24_r2 & !din_ready_3_24)begin
//       $display("overflow din_3_24");
//       $finish;
//   end
//    
//   if (din_almost_full_3_25) begin
//       $display("din_almost_full_3_25");
//   end  
//   if (din_valid_3_25_r2 & !din_ready_3_25)begin
//       $display("overflow din_3_25");
//       $finish;
//   end
//    
//   if (din_almost_full_3_26) begin
//       $display("din_almost_full_3_26");
//   end  
//   if (din_valid_3_26_r2 & !din_ready_3_26)begin
//       $display("overflow din_3_26");
//       $finish;
//   end
//    
//   if (din_almost_full_3_27) begin
//       $display("din_almost_full_3_27");
//   end  
//   if (din_valid_3_27_r2 & !din_ready_3_27)begin
//       $display("overflow din_3_27");
//       $finish;
//   end
//    
//   if (din_almost_full_3_28) begin
//       $display("din_almost_full_3_28");
//   end  
//   if (din_valid_3_28_r2 & !din_ready_3_28)begin
//       $display("overflow din_3_28");
//       $finish;
//   end
//    
//   if (din_almost_full_3_29) begin
//       $display("din_almost_full_3_29");
//   end  
//   if (din_valid_3_29_r2 & !din_ready_3_29)begin
//       $display("overflow din_3_29");
//       $finish;
//   end
//    
//   if (din_almost_full_3_30) begin
//       $display("din_almost_full_3_30");
//   end  
//   if (din_valid_3_30_r2 & !din_ready_3_30)begin
//       $display("overflow din_3_30");
//       $finish;
//   end
//    
//   if (din_almost_full_3_31) begin
//       $display("din_almost_full_3_31");
//   end  
//   if (din_valid_3_31_r2 & !din_ready_3_31)begin
//       $display("overflow din_3_31");
//       $finish;
//   end
//    
//    
//    
//   if (din_almost_full_4_0) begin
//       $display("din_almost_full_4_0");
//   end  
//   if (din_valid_4_0_r2 & !din_ready_4_0)begin
//       $display("overflow din_4_0");
//       $finish;
//   end
//    
//   if (din_almost_full_4_1) begin
//       $display("din_almost_full_4_1");
//   end  
//   if (din_valid_4_1_r2 & !din_ready_4_1)begin
//       $display("overflow din_4_1");
//       $finish;
//   end
//    
//   if (din_almost_full_4_2) begin
//       $display("din_almost_full_4_2");
//   end  
//   if (din_valid_4_2_r2 & !din_ready_4_2)begin
//       $display("overflow din_4_2");
//       $finish;
//   end
//    
//   if (din_almost_full_4_3) begin
//       $display("din_almost_full_4_3");
//   end  
//   if (din_valid_4_3_r2 & !din_ready_4_3)begin
//       $display("overflow din_4_3");
//       $finish;
//   end
//    
//   if (din_almost_full_4_4) begin
//       $display("din_almost_full_4_4");
//   end  
//   if (din_valid_4_4_r2 & !din_ready_4_4)begin
//       $display("overflow din_4_4");
//       $finish;
//   end
//    
//   if (din_almost_full_4_5) begin
//       $display("din_almost_full_4_5");
//   end  
//   if (din_valid_4_5_r2 & !din_ready_4_5)begin
//       $display("overflow din_4_5");
//       $finish;
//   end
//    
//   if (din_almost_full_4_6) begin
//       $display("din_almost_full_4_6");
//   end  
//   if (din_valid_4_6_r2 & !din_ready_4_6)begin
//       $display("overflow din_4_6");
//       $finish;
//   end
//    
//   if (din_almost_full_4_7) begin
//       $display("din_almost_full_4_7");
//   end  
//   if (din_valid_4_7_r2 & !din_ready_4_7)begin
//       $display("overflow din_4_7");
//       $finish;
//   end
//    
//   if (din_almost_full_4_8) begin
//       $display("din_almost_full_4_8");
//   end  
//   if (din_valid_4_8_r2 & !din_ready_4_8)begin
//       $display("overflow din_4_8");
//       $finish;
//   end
//    
//   if (din_almost_full_4_9) begin
//       $display("din_almost_full_4_9");
//   end  
//   if (din_valid_4_9_r2 & !din_ready_4_9)begin
//       $display("overflow din_4_9");
//       $finish;
//   end
//    
//   if (din_almost_full_4_10) begin
//       $display("din_almost_full_4_10");
//   end  
//   if (din_valid_4_10_r2 & !din_ready_4_10)begin
//       $display("overflow din_4_10");
//       $finish;
//   end
//    
//   if (din_almost_full_4_11) begin
//       $display("din_almost_full_4_11");
//   end  
//   if (din_valid_4_11_r2 & !din_ready_4_11)begin
//       $display("overflow din_4_11");
//       $finish;
//   end
//    
//   if (din_almost_full_4_12) begin
//       $display("din_almost_full_4_12");
//   end  
//   if (din_valid_4_12_r2 & !din_ready_4_12)begin
//       $display("overflow din_4_12");
//       $finish;
//   end
//    
//   if (din_almost_full_4_13) begin
//       $display("din_almost_full_4_13");
//   end  
//   if (din_valid_4_13_r2 & !din_ready_4_13)begin
//       $display("overflow din_4_13");
//       $finish;
//   end
//    
//   if (din_almost_full_4_14) begin
//       $display("din_almost_full_4_14");
//   end  
//   if (din_valid_4_14_r2 & !din_ready_4_14)begin
//       $display("overflow din_4_14");
//       $finish;
//   end
//    
//   if (din_almost_full_4_15) begin
//       $display("din_almost_full_4_15");
//   end  
//   if (din_valid_4_15_r2 & !din_ready_4_15)begin
//       $display("overflow din_4_15");
//       $finish;
//   end
//    
//   if (din_almost_full_4_16) begin
//       $display("din_almost_full_4_16");
//   end  
//   if (din_valid_4_16_r2 & !din_ready_4_16)begin
//       $display("overflow din_4_16");
//       $finish;
//   end
//    
//   if (din_almost_full_4_17) begin
//       $display("din_almost_full_4_17");
//   end  
//   if (din_valid_4_17_r2 & !din_ready_4_17)begin
//       $display("overflow din_4_17");
//       $finish;
//   end
//    
//   if (din_almost_full_4_18) begin
//       $display("din_almost_full_4_18");
//   end  
//   if (din_valid_4_18_r2 & !din_ready_4_18)begin
//       $display("overflow din_4_18");
//       $finish;
//   end
//    
//   if (din_almost_full_4_19) begin
//       $display("din_almost_full_4_19");
//   end  
//   if (din_valid_4_19_r2 & !din_ready_4_19)begin
//       $display("overflow din_4_19");
//       $finish;
//   end
//    
//   if (din_almost_full_4_20) begin
//       $display("din_almost_full_4_20");
//   end  
//   if (din_valid_4_20_r2 & !din_ready_4_20)begin
//       $display("overflow din_4_20");
//       $finish;
//   end
//    
//   if (din_almost_full_4_21) begin
//       $display("din_almost_full_4_21");
//   end  
//   if (din_valid_4_21_r2 & !din_ready_4_21)begin
//       $display("overflow din_4_21");
//       $finish;
//   end
//    
//   if (din_almost_full_4_22) begin
//       $display("din_almost_full_4_22");
//   end  
//   if (din_valid_4_22_r2 & !din_ready_4_22)begin
//       $display("overflow din_4_22");
//       $finish;
//   end
//    
//   if (din_almost_full_4_23) begin
//       $display("din_almost_full_4_23");
//   end  
//   if (din_valid_4_23_r2 & !din_ready_4_23)begin
//       $display("overflow din_4_23");
//       $finish;
//   end
//    
//   if (din_almost_full_4_24) begin
//       $display("din_almost_full_4_24");
//   end  
//   if (din_valid_4_24_r2 & !din_ready_4_24)begin
//       $display("overflow din_4_24");
//       $finish;
//   end
//    
//   if (din_almost_full_4_25) begin
//       $display("din_almost_full_4_25");
//   end  
//   if (din_valid_4_25_r2 & !din_ready_4_25)begin
//       $display("overflow din_4_25");
//       $finish;
//   end
//    
//   if (din_almost_full_4_26) begin
//       $display("din_almost_full_4_26");
//   end  
//   if (din_valid_4_26_r2 & !din_ready_4_26)begin
//       $display("overflow din_4_26");
//       $finish;
//   end
//    
//   if (din_almost_full_4_27) begin
//       $display("din_almost_full_4_27");
//   end  
//   if (din_valid_4_27_r2 & !din_ready_4_27)begin
//       $display("overflow din_4_27");
//       $finish;
//   end
//    
//   if (din_almost_full_4_28) begin
//       $display("din_almost_full_4_28");
//   end  
//   if (din_valid_4_28_r2 & !din_ready_4_28)begin
//       $display("overflow din_4_28");
//       $finish;
//   end
//    
//   if (din_almost_full_4_29) begin
//       $display("din_almost_full_4_29");
//   end  
//   if (din_valid_4_29_r2 & !din_ready_4_29)begin
//       $display("overflow din_4_29");
//       $finish;
//   end
//    
//   if (din_almost_full_4_30) begin
//       $display("din_almost_full_4_30");
//   end  
//   if (din_valid_4_30_r2 & !din_ready_4_30)begin
//       $display("overflow din_4_30");
//       $finish;
//   end
//    
//   if (din_almost_full_4_31) begin
//       $display("din_almost_full_4_31");
//   end  
//   if (din_valid_4_31_r2 & !din_ready_4_31)begin
//       $display("overflow din_4_31");
//       $finish;
//   end
//    
//    
//    
//   if (din_almost_full_5_0) begin
//       $display("din_almost_full_5_0");
//   end  
//   if (din_valid_5_0_r2 & !din_ready_5_0)begin
//       $display("overflow din_5_0");
//       $finish;
//   end
//    
//   if (din_almost_full_5_1) begin
//       $display("din_almost_full_5_1");
//   end  
//   if (din_valid_5_1_r2 & !din_ready_5_1)begin
//       $display("overflow din_5_1");
//       $finish;
//   end
//    
//   if (din_almost_full_5_2) begin
//       $display("din_almost_full_5_2");
//   end  
//   if (din_valid_5_2_r2 & !din_ready_5_2)begin
//       $display("overflow din_5_2");
//       $finish;
//   end
//    
//   if (din_almost_full_5_3) begin
//       $display("din_almost_full_5_3");
//   end  
//   if (din_valid_5_3_r2 & !din_ready_5_3)begin
//       $display("overflow din_5_3");
//       $finish;
//   end
//    
//   if (din_almost_full_5_4) begin
//       $display("din_almost_full_5_4");
//   end  
//   if (din_valid_5_4_r2 & !din_ready_5_4)begin
//       $display("overflow din_5_4");
//       $finish;
//   end
//    
//   if (din_almost_full_5_5) begin
//       $display("din_almost_full_5_5");
//   end  
//   if (din_valid_5_5_r2 & !din_ready_5_5)begin
//       $display("overflow din_5_5");
//       $finish;
//   end
//    
//   if (din_almost_full_5_6) begin
//       $display("din_almost_full_5_6");
//   end  
//   if (din_valid_5_6_r2 & !din_ready_5_6)begin
//       $display("overflow din_5_6");
//       $finish;
//   end
//    
//   if (din_almost_full_5_7) begin
//       $display("din_almost_full_5_7");
//   end  
//   if (din_valid_5_7_r2 & !din_ready_5_7)begin
//       $display("overflow din_5_7");
//       $finish;
//   end
//    
//   if (din_almost_full_5_8) begin
//       $display("din_almost_full_5_8");
//   end  
//   if (din_valid_5_8_r2 & !din_ready_5_8)begin
//       $display("overflow din_5_8");
//       $finish;
//   end
//    
//   if (din_almost_full_5_9) begin
//       $display("din_almost_full_5_9");
//   end  
//   if (din_valid_5_9_r2 & !din_ready_5_9)begin
//       $display("overflow din_5_9");
//       $finish;
//   end
//    
//   if (din_almost_full_5_10) begin
//       $display("din_almost_full_5_10");
//   end  
//   if (din_valid_5_10_r2 & !din_ready_5_10)begin
//       $display("overflow din_5_10");
//       $finish;
//   end
//    
//   if (din_almost_full_5_11) begin
//       $display("din_almost_full_5_11");
//   end  
//   if (din_valid_5_11_r2 & !din_ready_5_11)begin
//       $display("overflow din_5_11");
//       $finish;
//   end
//    
//   if (din_almost_full_5_12) begin
//       $display("din_almost_full_5_12");
//   end  
//   if (din_valid_5_12_r2 & !din_ready_5_12)begin
//       $display("overflow din_5_12");
//       $finish;
//   end
//    
//   if (din_almost_full_5_13) begin
//       $display("din_almost_full_5_13");
//   end  
//   if (din_valid_5_13_r2 & !din_ready_5_13)begin
//       $display("overflow din_5_13");
//       $finish;
//   end
//    
//   if (din_almost_full_5_14) begin
//       $display("din_almost_full_5_14");
//   end  
//   if (din_valid_5_14_r2 & !din_ready_5_14)begin
//       $display("overflow din_5_14");
//       $finish;
//   end
//    
//   if (din_almost_full_5_15) begin
//       $display("din_almost_full_5_15");
//   end  
//   if (din_valid_5_15_r2 & !din_ready_5_15)begin
//       $display("overflow din_5_15");
//       $finish;
//   end
//    
//   if (din_almost_full_5_16) begin
//       $display("din_almost_full_5_16");
//   end  
//   if (din_valid_5_16_r2 & !din_ready_5_16)begin
//       $display("overflow din_5_16");
//       $finish;
//   end
//    
//   if (din_almost_full_5_17) begin
//       $display("din_almost_full_5_17");
//   end  
//   if (din_valid_5_17_r2 & !din_ready_5_17)begin
//       $display("overflow din_5_17");
//       $finish;
//   end
//    
//   if (din_almost_full_5_18) begin
//       $display("din_almost_full_5_18");
//   end  
//   if (din_valid_5_18_r2 & !din_ready_5_18)begin
//       $display("overflow din_5_18");
//       $finish;
//   end
//    
//   if (din_almost_full_5_19) begin
//       $display("din_almost_full_5_19");
//   end  
//   if (din_valid_5_19_r2 & !din_ready_5_19)begin
//       $display("overflow din_5_19");
//       $finish;
//   end
//    
//   if (din_almost_full_5_20) begin
//       $display("din_almost_full_5_20");
//   end  
//   if (din_valid_5_20_r2 & !din_ready_5_20)begin
//       $display("overflow din_5_20");
//       $finish;
//   end
//    
//   if (din_almost_full_5_21) begin
//       $display("din_almost_full_5_21");
//   end  
//   if (din_valid_5_21_r2 & !din_ready_5_21)begin
//       $display("overflow din_5_21");
//       $finish;
//   end
//    
//   if (din_almost_full_5_22) begin
//       $display("din_almost_full_5_22");
//   end  
//   if (din_valid_5_22_r2 & !din_ready_5_22)begin
//       $display("overflow din_5_22");
//       $finish;
//   end
//    
//   if (din_almost_full_5_23) begin
//       $display("din_almost_full_5_23");
//   end  
//   if (din_valid_5_23_r2 & !din_ready_5_23)begin
//       $display("overflow din_5_23");
//       $finish;
//   end
//    
//   if (din_almost_full_5_24) begin
//       $display("din_almost_full_5_24");
//   end  
//   if (din_valid_5_24_r2 & !din_ready_5_24)begin
//       $display("overflow din_5_24");
//       $finish;
//   end
//    
//   if (din_almost_full_5_25) begin
//       $display("din_almost_full_5_25");
//   end  
//   if (din_valid_5_25_r2 & !din_ready_5_25)begin
//       $display("overflow din_5_25");
//       $finish;
//   end
//    
//   if (din_almost_full_5_26) begin
//       $display("din_almost_full_5_26");
//   end  
//   if (din_valid_5_26_r2 & !din_ready_5_26)begin
//       $display("overflow din_5_26");
//       $finish;
//   end
//    
//   if (din_almost_full_5_27) begin
//       $display("din_almost_full_5_27");
//   end  
//   if (din_valid_5_27_r2 & !din_ready_5_27)begin
//       $display("overflow din_5_27");
//       $finish;
//   end
//    
//   if (din_almost_full_5_28) begin
//       $display("din_almost_full_5_28");
//   end  
//   if (din_valid_5_28_r2 & !din_ready_5_28)begin
//       $display("overflow din_5_28");
//       $finish;
//   end
//    
//   if (din_almost_full_5_29) begin
//       $display("din_almost_full_5_29");
//   end  
//   if (din_valid_5_29_r2 & !din_ready_5_29)begin
//       $display("overflow din_5_29");
//       $finish;
//   end
//    
//   if (din_almost_full_5_30) begin
//       $display("din_almost_full_5_30");
//   end  
//   if (din_valid_5_30_r2 & !din_ready_5_30)begin
//       $display("overflow din_5_30");
//       $finish;
//   end
//    
//   if (din_almost_full_5_31) begin
//       $display("din_almost_full_5_31");
//   end  
//   if (din_valid_5_31_r2 & !din_ready_5_31)begin
//       $display("overflow din_5_31");
//       $finish;
//   end
//    
//    
//    
//   if (din_almost_full_6_0) begin
//       $display("din_almost_full_6_0");
//   end  
//   if (din_valid_6_0_r2 & !din_ready_6_0)begin
//       $display("overflow din_6_0");
//       $finish;
//   end
//    
//   if (din_almost_full_6_1) begin
//       $display("din_almost_full_6_1");
//   end  
//   if (din_valid_6_1_r2 & !din_ready_6_1)begin
//       $display("overflow din_6_1");
//       $finish;
//   end
//    
//   if (din_almost_full_6_2) begin
//       $display("din_almost_full_6_2");
//   end  
//   if (din_valid_6_2_r2 & !din_ready_6_2)begin
//       $display("overflow din_6_2");
//       $finish;
//   end
//    
//   if (din_almost_full_6_3) begin
//       $display("din_almost_full_6_3");
//   end  
//   if (din_valid_6_3_r2 & !din_ready_6_3)begin
//       $display("overflow din_6_3");
//       $finish;
//   end
//    
//   if (din_almost_full_6_4) begin
//       $display("din_almost_full_6_4");
//   end  
//   if (din_valid_6_4_r2 & !din_ready_6_4)begin
//       $display("overflow din_6_4");
//       $finish;
//   end
//    
//   if (din_almost_full_6_5) begin
//       $display("din_almost_full_6_5");
//   end  
//   if (din_valid_6_5_r2 & !din_ready_6_5)begin
//       $display("overflow din_6_5");
//       $finish;
//   end
//    
//   if (din_almost_full_6_6) begin
//       $display("din_almost_full_6_6");
//   end  
//   if (din_valid_6_6_r2 & !din_ready_6_6)begin
//       $display("overflow din_6_6");
//       $finish;
//   end
//    
//   if (din_almost_full_6_7) begin
//       $display("din_almost_full_6_7");
//   end  
//   if (din_valid_6_7_r2 & !din_ready_6_7)begin
//       $display("overflow din_6_7");
//       $finish;
//   end
//    
//   if (din_almost_full_6_8) begin
//       $display("din_almost_full_6_8");
//   end  
//   if (din_valid_6_8_r2 & !din_ready_6_8)begin
//       $display("overflow din_6_8");
//       $finish;
//   end
//    
//   if (din_almost_full_6_9) begin
//       $display("din_almost_full_6_9");
//   end  
//   if (din_valid_6_9_r2 & !din_ready_6_9)begin
//       $display("overflow din_6_9");
//       $finish;
//   end
//    
//   if (din_almost_full_6_10) begin
//       $display("din_almost_full_6_10");
//   end  
//   if (din_valid_6_10_r2 & !din_ready_6_10)begin
//       $display("overflow din_6_10");
//       $finish;
//   end
//    
//   if (din_almost_full_6_11) begin
//       $display("din_almost_full_6_11");
//   end  
//   if (din_valid_6_11_r2 & !din_ready_6_11)begin
//       $display("overflow din_6_11");
//       $finish;
//   end
//    
//   if (din_almost_full_6_12) begin
//       $display("din_almost_full_6_12");
//   end  
//   if (din_valid_6_12_r2 & !din_ready_6_12)begin
//       $display("overflow din_6_12");
//       $finish;
//   end
//    
//   if (din_almost_full_6_13) begin
//       $display("din_almost_full_6_13");
//   end  
//   if (din_valid_6_13_r2 & !din_ready_6_13)begin
//       $display("overflow din_6_13");
//       $finish;
//   end
//    
//   if (din_almost_full_6_14) begin
//       $display("din_almost_full_6_14");
//   end  
//   if (din_valid_6_14_r2 & !din_ready_6_14)begin
//       $display("overflow din_6_14");
//       $finish;
//   end
//    
//   if (din_almost_full_6_15) begin
//       $display("din_almost_full_6_15");
//   end  
//   if (din_valid_6_15_r2 & !din_ready_6_15)begin
//       $display("overflow din_6_15");
//       $finish;
//   end
//    
//   if (din_almost_full_6_16) begin
//       $display("din_almost_full_6_16");
//   end  
//   if (din_valid_6_16_r2 & !din_ready_6_16)begin
//       $display("overflow din_6_16");
//       $finish;
//   end
//    
//   if (din_almost_full_6_17) begin
//       $display("din_almost_full_6_17");
//   end  
//   if (din_valid_6_17_r2 & !din_ready_6_17)begin
//       $display("overflow din_6_17");
//       $finish;
//   end
//    
//   if (din_almost_full_6_18) begin
//       $display("din_almost_full_6_18");
//   end  
//   if (din_valid_6_18_r2 & !din_ready_6_18)begin
//       $display("overflow din_6_18");
//       $finish;
//   end
//    
//   if (din_almost_full_6_19) begin
//       $display("din_almost_full_6_19");
//   end  
//   if (din_valid_6_19_r2 & !din_ready_6_19)begin
//       $display("overflow din_6_19");
//       $finish;
//   end
//    
//   if (din_almost_full_6_20) begin
//       $display("din_almost_full_6_20");
//   end  
//   if (din_valid_6_20_r2 & !din_ready_6_20)begin
//       $display("overflow din_6_20");
//       $finish;
//   end
//    
//   if (din_almost_full_6_21) begin
//       $display("din_almost_full_6_21");
//   end  
//   if (din_valid_6_21_r2 & !din_ready_6_21)begin
//       $display("overflow din_6_21");
//       $finish;
//   end
//    
//   if (din_almost_full_6_22) begin
//       $display("din_almost_full_6_22");
//   end  
//   if (din_valid_6_22_r2 & !din_ready_6_22)begin
//       $display("overflow din_6_22");
//       $finish;
//   end
//    
//   if (din_almost_full_6_23) begin
//       $display("din_almost_full_6_23");
//   end  
//   if (din_valid_6_23_r2 & !din_ready_6_23)begin
//       $display("overflow din_6_23");
//       $finish;
//   end
//    
//   if (din_almost_full_6_24) begin
//       $display("din_almost_full_6_24");
//   end  
//   if (din_valid_6_24_r2 & !din_ready_6_24)begin
//       $display("overflow din_6_24");
//       $finish;
//   end
//    
//   if (din_almost_full_6_25) begin
//       $display("din_almost_full_6_25");
//   end  
//   if (din_valid_6_25_r2 & !din_ready_6_25)begin
//       $display("overflow din_6_25");
//       $finish;
//   end
//    
//   if (din_almost_full_6_26) begin
//       $display("din_almost_full_6_26");
//   end  
//   if (din_valid_6_26_r2 & !din_ready_6_26)begin
//       $display("overflow din_6_26");
//       $finish;
//   end
//    
//   if (din_almost_full_6_27) begin
//       $display("din_almost_full_6_27");
//   end  
//   if (din_valid_6_27_r2 & !din_ready_6_27)begin
//       $display("overflow din_6_27");
//       $finish;
//   end
//    
//   if (din_almost_full_6_28) begin
//       $display("din_almost_full_6_28");
//   end  
//   if (din_valid_6_28_r2 & !din_ready_6_28)begin
//       $display("overflow din_6_28");
//       $finish;
//   end
//    
//   if (din_almost_full_6_29) begin
//       $display("din_almost_full_6_29");
//   end  
//   if (din_valid_6_29_r2 & !din_ready_6_29)begin
//       $display("overflow din_6_29");
//       $finish;
//   end
//    
//   if (din_almost_full_6_30) begin
//       $display("din_almost_full_6_30");
//   end  
//   if (din_valid_6_30_r2 & !din_ready_6_30)begin
//       $display("overflow din_6_30");
//       $finish;
//   end
//    
//   if (din_almost_full_6_31) begin
//       $display("din_almost_full_6_31");
//   end  
//   if (din_valid_6_31_r2 & !din_ready_6_31)begin
//       $display("overflow din_6_31");
//       $finish;
//   end
//    
//    
//    
//   if (din_almost_full_7_0) begin
//       $display("din_almost_full_7_0");
//   end  
//   if (din_valid_7_0_r2 & !din_ready_7_0)begin
//       $display("overflow din_7_0");
//       $finish;
//   end
//    
//   if (din_almost_full_7_1) begin
//       $display("din_almost_full_7_1");
//   end  
//   if (din_valid_7_1_r2 & !din_ready_7_1)begin
//       $display("overflow din_7_1");
//       $finish;
//   end
//    
//   if (din_almost_full_7_2) begin
//       $display("din_almost_full_7_2");
//   end  
//   if (din_valid_7_2_r2 & !din_ready_7_2)begin
//       $display("overflow din_7_2");
//       $finish;
//   end
//    
//   if (din_almost_full_7_3) begin
//       $display("din_almost_full_7_3");
//   end  
//   if (din_valid_7_3_r2 & !din_ready_7_3)begin
//       $display("overflow din_7_3");
//       $finish;
//   end
//    
//   if (din_almost_full_7_4) begin
//       $display("din_almost_full_7_4");
//   end  
//   if (din_valid_7_4_r2 & !din_ready_7_4)begin
//       $display("overflow din_7_4");
//       $finish;
//   end
//    
//   if (din_almost_full_7_5) begin
//       $display("din_almost_full_7_5");
//   end  
//   if (din_valid_7_5_r2 & !din_ready_7_5)begin
//       $display("overflow din_7_5");
//       $finish;
//   end
//    
//   if (din_almost_full_7_6) begin
//       $display("din_almost_full_7_6");
//   end  
//   if (din_valid_7_6_r2 & !din_ready_7_6)begin
//       $display("overflow din_7_6");
//       $finish;
//   end
//    
//   if (din_almost_full_7_7) begin
//       $display("din_almost_full_7_7");
//   end  
//   if (din_valid_7_7_r2 & !din_ready_7_7)begin
//       $display("overflow din_7_7");
//       $finish;
//   end
//    
//   if (din_almost_full_7_8) begin
//       $display("din_almost_full_7_8");
//   end  
//   if (din_valid_7_8_r2 & !din_ready_7_8)begin
//       $display("overflow din_7_8");
//       $finish;
//   end
//    
//   if (din_almost_full_7_9) begin
//       $display("din_almost_full_7_9");
//   end  
//   if (din_valid_7_9_r2 & !din_ready_7_9)begin
//       $display("overflow din_7_9");
//       $finish;
//   end
//    
//   if (din_almost_full_7_10) begin
//       $display("din_almost_full_7_10");
//   end  
//   if (din_valid_7_10_r2 & !din_ready_7_10)begin
//       $display("overflow din_7_10");
//       $finish;
//   end
//    
//   if (din_almost_full_7_11) begin
//       $display("din_almost_full_7_11");
//   end  
//   if (din_valid_7_11_r2 & !din_ready_7_11)begin
//       $display("overflow din_7_11");
//       $finish;
//   end
//    
//   if (din_almost_full_7_12) begin
//       $display("din_almost_full_7_12");
//   end  
//   if (din_valid_7_12_r2 & !din_ready_7_12)begin
//       $display("overflow din_7_12");
//       $finish;
//   end
//    
//   if (din_almost_full_7_13) begin
//       $display("din_almost_full_7_13");
//   end  
//   if (din_valid_7_13_r2 & !din_ready_7_13)begin
//       $display("overflow din_7_13");
//       $finish;
//   end
//    
//   if (din_almost_full_7_14) begin
//       $display("din_almost_full_7_14");
//   end  
//   if (din_valid_7_14_r2 & !din_ready_7_14)begin
//       $display("overflow din_7_14");
//       $finish;
//   end
//    
//   if (din_almost_full_7_15) begin
//       $display("din_almost_full_7_15");
//   end  
//   if (din_valid_7_15_r2 & !din_ready_7_15)begin
//       $display("overflow din_7_15");
//       $finish;
//   end
//    
//   if (din_almost_full_7_16) begin
//       $display("din_almost_full_7_16");
//   end  
//   if (din_valid_7_16_r2 & !din_ready_7_16)begin
//       $display("overflow din_7_16");
//       $finish;
//   end
//    
//   if (din_almost_full_7_17) begin
//       $display("din_almost_full_7_17");
//   end  
//   if (din_valid_7_17_r2 & !din_ready_7_17)begin
//       $display("overflow din_7_17");
//       $finish;
//   end
//    
//   if (din_almost_full_7_18) begin
//       $display("din_almost_full_7_18");
//   end  
//   if (din_valid_7_18_r2 & !din_ready_7_18)begin
//       $display("overflow din_7_18");
//       $finish;
//   end
//    
//   if (din_almost_full_7_19) begin
//       $display("din_almost_full_7_19");
//   end  
//   if (din_valid_7_19_r2 & !din_ready_7_19)begin
//       $display("overflow din_7_19");
//       $finish;
//   end
//    
//   if (din_almost_full_7_20) begin
//       $display("din_almost_full_7_20");
//   end  
//   if (din_valid_7_20_r2 & !din_ready_7_20)begin
//       $display("overflow din_7_20");
//       $finish;
//   end
//    
//   if (din_almost_full_7_21) begin
//       $display("din_almost_full_7_21");
//   end  
//   if (din_valid_7_21_r2 & !din_ready_7_21)begin
//       $display("overflow din_7_21");
//       $finish;
//   end
//    
//   if (din_almost_full_7_22) begin
//       $display("din_almost_full_7_22");
//   end  
//   if (din_valid_7_22_r2 & !din_ready_7_22)begin
//       $display("overflow din_7_22");
//       $finish;
//   end
//    
//   if (din_almost_full_7_23) begin
//       $display("din_almost_full_7_23");
//   end  
//   if (din_valid_7_23_r2 & !din_ready_7_23)begin
//       $display("overflow din_7_23");
//       $finish;
//   end
//    
//   if (din_almost_full_7_24) begin
//       $display("din_almost_full_7_24");
//   end  
//   if (din_valid_7_24_r2 & !din_ready_7_24)begin
//       $display("overflow din_7_24");
//       $finish;
//   end
//    
//   if (din_almost_full_7_25) begin
//       $display("din_almost_full_7_25");
//   end  
//   if (din_valid_7_25_r2 & !din_ready_7_25)begin
//       $display("overflow din_7_25");
//       $finish;
//   end
//    
//   if (din_almost_full_7_26) begin
//       $display("din_almost_full_7_26");
//   end  
//   if (din_valid_7_26_r2 & !din_ready_7_26)begin
//       $display("overflow din_7_26");
//       $finish;
//   end
//    
//   if (din_almost_full_7_27) begin
//       $display("din_almost_full_7_27");
//   end  
//   if (din_valid_7_27_r2 & !din_ready_7_27)begin
//       $display("overflow din_7_27");
//       $finish;
//   end
//    
//   if (din_almost_full_7_28) begin
//       $display("din_almost_full_7_28");
//   end  
//   if (din_valid_7_28_r2 & !din_ready_7_28)begin
//       $display("overflow din_7_28");
//       $finish;
//   end
//    
//   if (din_almost_full_7_29) begin
//       $display("din_almost_full_7_29");
//   end  
//   if (din_valid_7_29_r2 & !din_ready_7_29)begin
//       $display("overflow din_7_29");
//       $finish;
//   end
//    
//   if (din_almost_full_7_30) begin
//       $display("din_almost_full_7_30");
//   end  
//   if (din_valid_7_30_r2 & !din_ready_7_30)begin
//       $display("overflow din_7_30");
//       $finish;
//   end
//    
//   if (din_almost_full_7_31) begin
//       $display("din_almost_full_7_31");
//   end  
//   if (din_valid_7_31_r2 & !din_ready_7_31)begin
//       $display("overflow din_7_31");
//       $finish;
//   end
//    
//   //end

always @ (posedge front_clk) begin
    if(front_rst)begin
        in_pkt_cnt <= 0;
    end else begin
        if (in_pkt_valid & in_pkt_eop & in_pkt_ready) begin
            in_pkt_cnt <= in_pkt_cnt + 1;
        end
    end
end

always @ (posedge back_clk) begin
    if(back_rst)begin
        out_rule_cnt <= 0;
        out_rule_last_cnt <= 0;
    end else begin
        if(out_usr_valid & out_usr_ready)begin
            out_rule_cnt <= out_rule_cnt + 1;
            if(out_usr_eop)begin
                out_rule_last_cnt <= out_rule_last_cnt + 1;
            end
        end
    end
end


always@(posedge front_clk)begin
    din_valid_0_0 <= out_new_pkt | hash_out_valid_filter_0_0;
    din_valid_0_0_r1 <= din_valid_0_0;
    din_valid_0_0_r2 <= din_valid_0_0_r1;

    din_0_0.data <= hash_out_valid_filter_0_0 ? hash_out_0_0 : 0;
    din_0_0.last <= out_new_pkt;
    din_0_0.bucket <= 0;


    din_0_0_r1 <= din_0_0;
    din_0_0_r2 <= din_0_0_r1;
    din_valid_0_1 <= out_new_pkt | hash_out_valid_filter_0_1;
    din_valid_0_1_r1 <= din_valid_0_1;
    din_valid_0_1_r2 <= din_valid_0_1_r1;

    din_0_1.data <= hash_out_valid_filter_0_1 ? hash_out_0_1 : 0;
    din_0_1.last <= out_new_pkt;
    din_0_1.bucket <= 0;


    din_0_1_r1 <= din_0_1;
    din_0_1_r2 <= din_0_1_r1;
    din_valid_0_2 <= out_new_pkt | hash_out_valid_filter_0_2;
    din_valid_0_2_r1 <= din_valid_0_2;
    din_valid_0_2_r2 <= din_valid_0_2_r1;

    din_0_2.data <= hash_out_valid_filter_0_2 ? hash_out_0_2 : 0;
    din_0_2.last <= out_new_pkt;
    din_0_2.bucket <= 0;


    din_0_2_r1 <= din_0_2;
    din_0_2_r2 <= din_0_2_r1;
    din_valid_0_3 <= out_new_pkt | hash_out_valid_filter_0_3;
    din_valid_0_3_r1 <= din_valid_0_3;
    din_valid_0_3_r2 <= din_valid_0_3_r1;

    din_0_3.data <= hash_out_valid_filter_0_3 ? hash_out_0_3 : 0;
    din_0_3.last <= out_new_pkt;
    din_0_3.bucket <= 0;


    din_0_3_r1 <= din_0_3;
    din_0_3_r2 <= din_0_3_r1;
    din_valid_0_4 <= out_new_pkt | hash_out_valid_filter_0_4;
    din_valid_0_4_r1 <= din_valid_0_4;
    din_valid_0_4_r2 <= din_valid_0_4_r1;

    din_0_4.data <= hash_out_valid_filter_0_4 ? hash_out_0_4 : 0;
    din_0_4.last <= out_new_pkt;
    din_0_4.bucket <= 0;


    din_0_4_r1 <= din_0_4;
    din_0_4_r2 <= din_0_4_r1;
    din_valid_0_5 <= out_new_pkt | hash_out_valid_filter_0_5;
    din_valid_0_5_r1 <= din_valid_0_5;
    din_valid_0_5_r2 <= din_valid_0_5_r1;

    din_0_5.data <= hash_out_valid_filter_0_5 ? hash_out_0_5 : 0;
    din_0_5.last <= out_new_pkt;
    din_0_5.bucket <= 0;


    din_0_5_r1 <= din_0_5;
    din_0_5_r2 <= din_0_5_r1;
    din_valid_0_6 <= out_new_pkt | hash_out_valid_filter_0_6;
    din_valid_0_6_r1 <= din_valid_0_6;
    din_valid_0_6_r2 <= din_valid_0_6_r1;

    din_0_6.data <= hash_out_valid_filter_0_6 ? hash_out_0_6 : 0;
    din_0_6.last <= out_new_pkt;
    din_0_6.bucket <= 0;


    din_0_6_r1 <= din_0_6;
    din_0_6_r2 <= din_0_6_r1;
    din_valid_0_7 <= out_new_pkt | hash_out_valid_filter_0_7;
    din_valid_0_7_r1 <= din_valid_0_7;
    din_valid_0_7_r2 <= din_valid_0_7_r1;

    din_0_7.data <= hash_out_valid_filter_0_7 ? hash_out_0_7 : 0;
    din_0_7.last <= out_new_pkt;
    din_0_7.bucket <= 0;


    din_0_7_r1 <= din_0_7;
    din_0_7_r2 <= din_0_7_r1;
    din_valid_0_8 <= out_new_pkt | hash_out_valid_filter_0_8;
    din_valid_0_8_r1 <= din_valid_0_8;
    din_valid_0_8_r2 <= din_valid_0_8_r1;

    din_0_8.data <= hash_out_valid_filter_0_8 ? hash_out_0_8 : 0;
    din_0_8.last <= out_new_pkt;
    din_0_8.bucket <= 0;


    din_0_8_r1 <= din_0_8;
    din_0_8_r2 <= din_0_8_r1;
    din_valid_0_9 <= out_new_pkt | hash_out_valid_filter_0_9;
    din_valid_0_9_r1 <= din_valid_0_9;
    din_valid_0_9_r2 <= din_valid_0_9_r1;

    din_0_9.data <= hash_out_valid_filter_0_9 ? hash_out_0_9 : 0;
    din_0_9.last <= out_new_pkt;
    din_0_9.bucket <= 0;


    din_0_9_r1 <= din_0_9;
    din_0_9_r2 <= din_0_9_r1;
    din_valid_0_10 <= out_new_pkt | hash_out_valid_filter_0_10;
    din_valid_0_10_r1 <= din_valid_0_10;
    din_valid_0_10_r2 <= din_valid_0_10_r1;

    din_0_10.data <= hash_out_valid_filter_0_10 ? hash_out_0_10 : 0;
    din_0_10.last <= out_new_pkt;
    din_0_10.bucket <= 0;


    din_0_10_r1 <= din_0_10;
    din_0_10_r2 <= din_0_10_r1;
    din_valid_0_11 <= out_new_pkt | hash_out_valid_filter_0_11;
    din_valid_0_11_r1 <= din_valid_0_11;
    din_valid_0_11_r2 <= din_valid_0_11_r1;

    din_0_11.data <= hash_out_valid_filter_0_11 ? hash_out_0_11 : 0;
    din_0_11.last <= out_new_pkt;
    din_0_11.bucket <= 0;


    din_0_11_r1 <= din_0_11;
    din_0_11_r2 <= din_0_11_r1;
    din_valid_0_12 <= out_new_pkt | hash_out_valid_filter_0_12;
    din_valid_0_12_r1 <= din_valid_0_12;
    din_valid_0_12_r2 <= din_valid_0_12_r1;

    din_0_12.data <= hash_out_valid_filter_0_12 ? hash_out_0_12 : 0;
    din_0_12.last <= out_new_pkt;
    din_0_12.bucket <= 0;


    din_0_12_r1 <= din_0_12;
    din_0_12_r2 <= din_0_12_r1;
    din_valid_0_13 <= out_new_pkt | hash_out_valid_filter_0_13;
    din_valid_0_13_r1 <= din_valid_0_13;
    din_valid_0_13_r2 <= din_valid_0_13_r1;

    din_0_13.data <= hash_out_valid_filter_0_13 ? hash_out_0_13 : 0;
    din_0_13.last <= out_new_pkt;
    din_0_13.bucket <= 0;


    din_0_13_r1 <= din_0_13;
    din_0_13_r2 <= din_0_13_r1;
    din_valid_0_14 <= out_new_pkt | hash_out_valid_filter_0_14;
    din_valid_0_14_r1 <= din_valid_0_14;
    din_valid_0_14_r2 <= din_valid_0_14_r1;

    din_0_14.data <= hash_out_valid_filter_0_14 ? hash_out_0_14 : 0;
    din_0_14.last <= out_new_pkt;
    din_0_14.bucket <= 0;


    din_0_14_r1 <= din_0_14;
    din_0_14_r2 <= din_0_14_r1;
    din_valid_0_15 <= out_new_pkt | hash_out_valid_filter_0_15;
    din_valid_0_15_r1 <= din_valid_0_15;
    din_valid_0_15_r2 <= din_valid_0_15_r1;

    din_0_15.data <= hash_out_valid_filter_0_15 ? hash_out_0_15 : 0;
    din_0_15.last <= out_new_pkt;
    din_0_15.bucket <= 0;


    din_0_15_r1 <= din_0_15;
    din_0_15_r2 <= din_0_15_r1;
    din_valid_0_16 <= out_new_pkt | hash_out_valid_filter_0_16;
    din_valid_0_16_r1 <= din_valid_0_16;
    din_valid_0_16_r2 <= din_valid_0_16_r1;

    din_0_16.data <= hash_out_valid_filter_0_16 ? hash_out_0_16 : 0;
    din_0_16.last <= out_new_pkt;
    din_0_16.bucket <= 0;


    din_0_16_r1 <= din_0_16;
    din_0_16_r2 <= din_0_16_r1;
    din_valid_0_17 <= out_new_pkt | hash_out_valid_filter_0_17;
    din_valid_0_17_r1 <= din_valid_0_17;
    din_valid_0_17_r2 <= din_valid_0_17_r1;

    din_0_17.data <= hash_out_valid_filter_0_17 ? hash_out_0_17 : 0;
    din_0_17.last <= out_new_pkt;
    din_0_17.bucket <= 0;


    din_0_17_r1 <= din_0_17;
    din_0_17_r2 <= din_0_17_r1;
    din_valid_0_18 <= out_new_pkt | hash_out_valid_filter_0_18;
    din_valid_0_18_r1 <= din_valid_0_18;
    din_valid_0_18_r2 <= din_valid_0_18_r1;

    din_0_18.data <= hash_out_valid_filter_0_18 ? hash_out_0_18 : 0;
    din_0_18.last <= out_new_pkt;
    din_0_18.bucket <= 0;


    din_0_18_r1 <= din_0_18;
    din_0_18_r2 <= din_0_18_r1;
    din_valid_0_19 <= out_new_pkt | hash_out_valid_filter_0_19;
    din_valid_0_19_r1 <= din_valid_0_19;
    din_valid_0_19_r2 <= din_valid_0_19_r1;

    din_0_19.data <= hash_out_valid_filter_0_19 ? hash_out_0_19 : 0;
    din_0_19.last <= out_new_pkt;
    din_0_19.bucket <= 0;


    din_0_19_r1 <= din_0_19;
    din_0_19_r2 <= din_0_19_r1;
    din_valid_0_20 <= out_new_pkt | hash_out_valid_filter_0_20;
    din_valid_0_20_r1 <= din_valid_0_20;
    din_valid_0_20_r2 <= din_valid_0_20_r1;

    din_0_20.data <= hash_out_valid_filter_0_20 ? hash_out_0_20 : 0;
    din_0_20.last <= out_new_pkt;
    din_0_20.bucket <= 0;


    din_0_20_r1 <= din_0_20;
    din_0_20_r2 <= din_0_20_r1;
    din_valid_0_21 <= out_new_pkt | hash_out_valid_filter_0_21;
    din_valid_0_21_r1 <= din_valid_0_21;
    din_valid_0_21_r2 <= din_valid_0_21_r1;

    din_0_21.data <= hash_out_valid_filter_0_21 ? hash_out_0_21 : 0;
    din_0_21.last <= out_new_pkt;
    din_0_21.bucket <= 0;


    din_0_21_r1 <= din_0_21;
    din_0_21_r2 <= din_0_21_r1;
    din_valid_0_22 <= out_new_pkt | hash_out_valid_filter_0_22;
    din_valid_0_22_r1 <= din_valid_0_22;
    din_valid_0_22_r2 <= din_valid_0_22_r1;

    din_0_22.data <= hash_out_valid_filter_0_22 ? hash_out_0_22 : 0;
    din_0_22.last <= out_new_pkt;
    din_0_22.bucket <= 0;


    din_0_22_r1 <= din_0_22;
    din_0_22_r2 <= din_0_22_r1;
    din_valid_0_23 <= out_new_pkt | hash_out_valid_filter_0_23;
    din_valid_0_23_r1 <= din_valid_0_23;
    din_valid_0_23_r2 <= din_valid_0_23_r1;

    din_0_23.data <= hash_out_valid_filter_0_23 ? hash_out_0_23 : 0;
    din_0_23.last <= out_new_pkt;
    din_0_23.bucket <= 0;


    din_0_23_r1 <= din_0_23;
    din_0_23_r2 <= din_0_23_r1;
    din_valid_0_24 <= out_new_pkt | hash_out_valid_filter_0_24;
    din_valid_0_24_r1 <= din_valid_0_24;
    din_valid_0_24_r2 <= din_valid_0_24_r1;

    din_0_24.data <= hash_out_valid_filter_0_24 ? hash_out_0_24 : 0;
    din_0_24.last <= out_new_pkt;
    din_0_24.bucket <= 0;


    din_0_24_r1 <= din_0_24;
    din_0_24_r2 <= din_0_24_r1;
    din_valid_0_25 <= out_new_pkt | hash_out_valid_filter_0_25;
    din_valid_0_25_r1 <= din_valid_0_25;
    din_valid_0_25_r2 <= din_valid_0_25_r1;

    din_0_25.data <= hash_out_valid_filter_0_25 ? hash_out_0_25 : 0;
    din_0_25.last <= out_new_pkt;
    din_0_25.bucket <= 0;


    din_0_25_r1 <= din_0_25;
    din_0_25_r2 <= din_0_25_r1;
    din_valid_0_26 <= out_new_pkt | hash_out_valid_filter_0_26;
    din_valid_0_26_r1 <= din_valid_0_26;
    din_valid_0_26_r2 <= din_valid_0_26_r1;

    din_0_26.data <= hash_out_valid_filter_0_26 ? hash_out_0_26 : 0;
    din_0_26.last <= out_new_pkt;
    din_0_26.bucket <= 0;


    din_0_26_r1 <= din_0_26;
    din_0_26_r2 <= din_0_26_r1;
    din_valid_0_27 <= out_new_pkt | hash_out_valid_filter_0_27;
    din_valid_0_27_r1 <= din_valid_0_27;
    din_valid_0_27_r2 <= din_valid_0_27_r1;

    din_0_27.data <= hash_out_valid_filter_0_27 ? hash_out_0_27 : 0;
    din_0_27.last <= out_new_pkt;
    din_0_27.bucket <= 0;


    din_0_27_r1 <= din_0_27;
    din_0_27_r2 <= din_0_27_r1;
    din_valid_0_28 <= out_new_pkt | hash_out_valid_filter_0_28;
    din_valid_0_28_r1 <= din_valid_0_28;
    din_valid_0_28_r2 <= din_valid_0_28_r1;

    din_0_28.data <= hash_out_valid_filter_0_28 ? hash_out_0_28 : 0;
    din_0_28.last <= out_new_pkt;
    din_0_28.bucket <= 0;


    din_0_28_r1 <= din_0_28;
    din_0_28_r2 <= din_0_28_r1;
    din_valid_0_29 <= out_new_pkt | hash_out_valid_filter_0_29;
    din_valid_0_29_r1 <= din_valid_0_29;
    din_valid_0_29_r2 <= din_valid_0_29_r1;

    din_0_29.data <= hash_out_valid_filter_0_29 ? hash_out_0_29 : 0;
    din_0_29.last <= out_new_pkt;
    din_0_29.bucket <= 0;


    din_0_29_r1 <= din_0_29;
    din_0_29_r2 <= din_0_29_r1;
    din_valid_0_30 <= out_new_pkt | hash_out_valid_filter_0_30;
    din_valid_0_30_r1 <= din_valid_0_30;
    din_valid_0_30_r2 <= din_valid_0_30_r1;

    din_0_30.data <= hash_out_valid_filter_0_30 ? hash_out_0_30 : 0;
    din_0_30.last <= out_new_pkt;
    din_0_30.bucket <= 0;


    din_0_30_r1 <= din_0_30;
    din_0_30_r2 <= din_0_30_r1;
    din_valid_0_31 <= out_new_pkt | hash_out_valid_filter_0_31;
    din_valid_0_31_r1 <= din_valid_0_31;
    din_valid_0_31_r2 <= din_valid_0_31_r1;

    din_0_31.data <= hash_out_valid_filter_0_31 ? hash_out_0_31 : 0;
    din_0_31.last <= out_new_pkt;
    din_0_31.bucket <= 0;


    din_0_31_r1 <= din_0_31;
    din_0_31_r2 <= din_0_31_r1;
    din_valid_1_0 <= out_new_pkt | hash_out_valid_filter_1_0;
    din_valid_1_0_r1 <= din_valid_1_0;
    din_valid_1_0_r2 <= din_valid_1_0_r1;

    din_1_0.data <= hash_out_valid_filter_1_0 ? hash_out_1_0 : 0;
    din_1_0.last <= out_new_pkt;
    din_1_0.bucket <= 1;


    din_1_0_r1 <= din_1_0;
    din_1_0_r2 <= din_1_0_r1;
    din_valid_1_1 <= out_new_pkt | hash_out_valid_filter_1_1;
    din_valid_1_1_r1 <= din_valid_1_1;
    din_valid_1_1_r2 <= din_valid_1_1_r1;

    din_1_1.data <= hash_out_valid_filter_1_1 ? hash_out_1_1 : 0;
    din_1_1.last <= out_new_pkt;
    din_1_1.bucket <= 1;


    din_1_1_r1 <= din_1_1;
    din_1_1_r2 <= din_1_1_r1;
    din_valid_1_2 <= out_new_pkt | hash_out_valid_filter_1_2;
    din_valid_1_2_r1 <= din_valid_1_2;
    din_valid_1_2_r2 <= din_valid_1_2_r1;

    din_1_2.data <= hash_out_valid_filter_1_2 ? hash_out_1_2 : 0;
    din_1_2.last <= out_new_pkt;
    din_1_2.bucket <= 1;


    din_1_2_r1 <= din_1_2;
    din_1_2_r2 <= din_1_2_r1;
    din_valid_1_3 <= out_new_pkt | hash_out_valid_filter_1_3;
    din_valid_1_3_r1 <= din_valid_1_3;
    din_valid_1_3_r2 <= din_valid_1_3_r1;

    din_1_3.data <= hash_out_valid_filter_1_3 ? hash_out_1_3 : 0;
    din_1_3.last <= out_new_pkt;
    din_1_3.bucket <= 1;


    din_1_3_r1 <= din_1_3;
    din_1_3_r2 <= din_1_3_r1;
    din_valid_1_4 <= out_new_pkt | hash_out_valid_filter_1_4;
    din_valid_1_4_r1 <= din_valid_1_4;
    din_valid_1_4_r2 <= din_valid_1_4_r1;

    din_1_4.data <= hash_out_valid_filter_1_4 ? hash_out_1_4 : 0;
    din_1_4.last <= out_new_pkt;
    din_1_4.bucket <= 1;


    din_1_4_r1 <= din_1_4;
    din_1_4_r2 <= din_1_4_r1;
    din_valid_1_5 <= out_new_pkt | hash_out_valid_filter_1_5;
    din_valid_1_5_r1 <= din_valid_1_5;
    din_valid_1_5_r2 <= din_valid_1_5_r1;

    din_1_5.data <= hash_out_valid_filter_1_5 ? hash_out_1_5 : 0;
    din_1_5.last <= out_new_pkt;
    din_1_5.bucket <= 1;


    din_1_5_r1 <= din_1_5;
    din_1_5_r2 <= din_1_5_r1;
    din_valid_1_6 <= out_new_pkt | hash_out_valid_filter_1_6;
    din_valid_1_6_r1 <= din_valid_1_6;
    din_valid_1_6_r2 <= din_valid_1_6_r1;

    din_1_6.data <= hash_out_valid_filter_1_6 ? hash_out_1_6 : 0;
    din_1_6.last <= out_new_pkt;
    din_1_6.bucket <= 1;


    din_1_6_r1 <= din_1_6;
    din_1_6_r2 <= din_1_6_r1;
    din_valid_1_7 <= out_new_pkt | hash_out_valid_filter_1_7;
    din_valid_1_7_r1 <= din_valid_1_7;
    din_valid_1_7_r2 <= din_valid_1_7_r1;

    din_1_7.data <= hash_out_valid_filter_1_7 ? hash_out_1_7 : 0;
    din_1_7.last <= out_new_pkt;
    din_1_7.bucket <= 1;


    din_1_7_r1 <= din_1_7;
    din_1_7_r2 <= din_1_7_r1;
    din_valid_1_8 <= out_new_pkt | hash_out_valid_filter_1_8;
    din_valid_1_8_r1 <= din_valid_1_8;
    din_valid_1_8_r2 <= din_valid_1_8_r1;

    din_1_8.data <= hash_out_valid_filter_1_8 ? hash_out_1_8 : 0;
    din_1_8.last <= out_new_pkt;
    din_1_8.bucket <= 1;


    din_1_8_r1 <= din_1_8;
    din_1_8_r2 <= din_1_8_r1;
    din_valid_1_9 <= out_new_pkt | hash_out_valid_filter_1_9;
    din_valid_1_9_r1 <= din_valid_1_9;
    din_valid_1_9_r2 <= din_valid_1_9_r1;

    din_1_9.data <= hash_out_valid_filter_1_9 ? hash_out_1_9 : 0;
    din_1_9.last <= out_new_pkt;
    din_1_9.bucket <= 1;


    din_1_9_r1 <= din_1_9;
    din_1_9_r2 <= din_1_9_r1;
    din_valid_1_10 <= out_new_pkt | hash_out_valid_filter_1_10;
    din_valid_1_10_r1 <= din_valid_1_10;
    din_valid_1_10_r2 <= din_valid_1_10_r1;

    din_1_10.data <= hash_out_valid_filter_1_10 ? hash_out_1_10 : 0;
    din_1_10.last <= out_new_pkt;
    din_1_10.bucket <= 1;


    din_1_10_r1 <= din_1_10;
    din_1_10_r2 <= din_1_10_r1;
    din_valid_1_11 <= out_new_pkt | hash_out_valid_filter_1_11;
    din_valid_1_11_r1 <= din_valid_1_11;
    din_valid_1_11_r2 <= din_valid_1_11_r1;

    din_1_11.data <= hash_out_valid_filter_1_11 ? hash_out_1_11 : 0;
    din_1_11.last <= out_new_pkt;
    din_1_11.bucket <= 1;


    din_1_11_r1 <= din_1_11;
    din_1_11_r2 <= din_1_11_r1;
    din_valid_1_12 <= out_new_pkt | hash_out_valid_filter_1_12;
    din_valid_1_12_r1 <= din_valid_1_12;
    din_valid_1_12_r2 <= din_valid_1_12_r1;

    din_1_12.data <= hash_out_valid_filter_1_12 ? hash_out_1_12 : 0;
    din_1_12.last <= out_new_pkt;
    din_1_12.bucket <= 1;


    din_1_12_r1 <= din_1_12;
    din_1_12_r2 <= din_1_12_r1;
    din_valid_1_13 <= out_new_pkt | hash_out_valid_filter_1_13;
    din_valid_1_13_r1 <= din_valid_1_13;
    din_valid_1_13_r2 <= din_valid_1_13_r1;

    din_1_13.data <= hash_out_valid_filter_1_13 ? hash_out_1_13 : 0;
    din_1_13.last <= out_new_pkt;
    din_1_13.bucket <= 1;


    din_1_13_r1 <= din_1_13;
    din_1_13_r2 <= din_1_13_r1;
    din_valid_1_14 <= out_new_pkt | hash_out_valid_filter_1_14;
    din_valid_1_14_r1 <= din_valid_1_14;
    din_valid_1_14_r2 <= din_valid_1_14_r1;

    din_1_14.data <= hash_out_valid_filter_1_14 ? hash_out_1_14 : 0;
    din_1_14.last <= out_new_pkt;
    din_1_14.bucket <= 1;


    din_1_14_r1 <= din_1_14;
    din_1_14_r2 <= din_1_14_r1;
    din_valid_1_15 <= out_new_pkt | hash_out_valid_filter_1_15;
    din_valid_1_15_r1 <= din_valid_1_15;
    din_valid_1_15_r2 <= din_valid_1_15_r1;

    din_1_15.data <= hash_out_valid_filter_1_15 ? hash_out_1_15 : 0;
    din_1_15.last <= out_new_pkt;
    din_1_15.bucket <= 1;


    din_1_15_r1 <= din_1_15;
    din_1_15_r2 <= din_1_15_r1;
    din_valid_1_16 <= out_new_pkt | hash_out_valid_filter_1_16;
    din_valid_1_16_r1 <= din_valid_1_16;
    din_valid_1_16_r2 <= din_valid_1_16_r1;

    din_1_16.data <= hash_out_valid_filter_1_16 ? hash_out_1_16 : 0;
    din_1_16.last <= out_new_pkt;
    din_1_16.bucket <= 1;


    din_1_16_r1 <= din_1_16;
    din_1_16_r2 <= din_1_16_r1;
    din_valid_1_17 <= out_new_pkt | hash_out_valid_filter_1_17;
    din_valid_1_17_r1 <= din_valid_1_17;
    din_valid_1_17_r2 <= din_valid_1_17_r1;

    din_1_17.data <= hash_out_valid_filter_1_17 ? hash_out_1_17 : 0;
    din_1_17.last <= out_new_pkt;
    din_1_17.bucket <= 1;


    din_1_17_r1 <= din_1_17;
    din_1_17_r2 <= din_1_17_r1;
    din_valid_1_18 <= out_new_pkt | hash_out_valid_filter_1_18;
    din_valid_1_18_r1 <= din_valid_1_18;
    din_valid_1_18_r2 <= din_valid_1_18_r1;

    din_1_18.data <= hash_out_valid_filter_1_18 ? hash_out_1_18 : 0;
    din_1_18.last <= out_new_pkt;
    din_1_18.bucket <= 1;


    din_1_18_r1 <= din_1_18;
    din_1_18_r2 <= din_1_18_r1;
    din_valid_1_19 <= out_new_pkt | hash_out_valid_filter_1_19;
    din_valid_1_19_r1 <= din_valid_1_19;
    din_valid_1_19_r2 <= din_valid_1_19_r1;

    din_1_19.data <= hash_out_valid_filter_1_19 ? hash_out_1_19 : 0;
    din_1_19.last <= out_new_pkt;
    din_1_19.bucket <= 1;


    din_1_19_r1 <= din_1_19;
    din_1_19_r2 <= din_1_19_r1;
    din_valid_1_20 <= out_new_pkt | hash_out_valid_filter_1_20;
    din_valid_1_20_r1 <= din_valid_1_20;
    din_valid_1_20_r2 <= din_valid_1_20_r1;

    din_1_20.data <= hash_out_valid_filter_1_20 ? hash_out_1_20 : 0;
    din_1_20.last <= out_new_pkt;
    din_1_20.bucket <= 1;


    din_1_20_r1 <= din_1_20;
    din_1_20_r2 <= din_1_20_r1;
    din_valid_1_21 <= out_new_pkt | hash_out_valid_filter_1_21;
    din_valid_1_21_r1 <= din_valid_1_21;
    din_valid_1_21_r2 <= din_valid_1_21_r1;

    din_1_21.data <= hash_out_valid_filter_1_21 ? hash_out_1_21 : 0;
    din_1_21.last <= out_new_pkt;
    din_1_21.bucket <= 1;


    din_1_21_r1 <= din_1_21;
    din_1_21_r2 <= din_1_21_r1;
    din_valid_1_22 <= out_new_pkt | hash_out_valid_filter_1_22;
    din_valid_1_22_r1 <= din_valid_1_22;
    din_valid_1_22_r2 <= din_valid_1_22_r1;

    din_1_22.data <= hash_out_valid_filter_1_22 ? hash_out_1_22 : 0;
    din_1_22.last <= out_new_pkt;
    din_1_22.bucket <= 1;


    din_1_22_r1 <= din_1_22;
    din_1_22_r2 <= din_1_22_r1;
    din_valid_1_23 <= out_new_pkt | hash_out_valid_filter_1_23;
    din_valid_1_23_r1 <= din_valid_1_23;
    din_valid_1_23_r2 <= din_valid_1_23_r1;

    din_1_23.data <= hash_out_valid_filter_1_23 ? hash_out_1_23 : 0;
    din_1_23.last <= out_new_pkt;
    din_1_23.bucket <= 1;


    din_1_23_r1 <= din_1_23;
    din_1_23_r2 <= din_1_23_r1;
    din_valid_1_24 <= out_new_pkt | hash_out_valid_filter_1_24;
    din_valid_1_24_r1 <= din_valid_1_24;
    din_valid_1_24_r2 <= din_valid_1_24_r1;

    din_1_24.data <= hash_out_valid_filter_1_24 ? hash_out_1_24 : 0;
    din_1_24.last <= out_new_pkt;
    din_1_24.bucket <= 1;


    din_1_24_r1 <= din_1_24;
    din_1_24_r2 <= din_1_24_r1;
    din_valid_1_25 <= out_new_pkt | hash_out_valid_filter_1_25;
    din_valid_1_25_r1 <= din_valid_1_25;
    din_valid_1_25_r2 <= din_valid_1_25_r1;

    din_1_25.data <= hash_out_valid_filter_1_25 ? hash_out_1_25 : 0;
    din_1_25.last <= out_new_pkt;
    din_1_25.bucket <= 1;


    din_1_25_r1 <= din_1_25;
    din_1_25_r2 <= din_1_25_r1;
    din_valid_1_26 <= out_new_pkt | hash_out_valid_filter_1_26;
    din_valid_1_26_r1 <= din_valid_1_26;
    din_valid_1_26_r2 <= din_valid_1_26_r1;

    din_1_26.data <= hash_out_valid_filter_1_26 ? hash_out_1_26 : 0;
    din_1_26.last <= out_new_pkt;
    din_1_26.bucket <= 1;


    din_1_26_r1 <= din_1_26;
    din_1_26_r2 <= din_1_26_r1;
    din_valid_1_27 <= out_new_pkt | hash_out_valid_filter_1_27;
    din_valid_1_27_r1 <= din_valid_1_27;
    din_valid_1_27_r2 <= din_valid_1_27_r1;

    din_1_27.data <= hash_out_valid_filter_1_27 ? hash_out_1_27 : 0;
    din_1_27.last <= out_new_pkt;
    din_1_27.bucket <= 1;


    din_1_27_r1 <= din_1_27;
    din_1_27_r2 <= din_1_27_r1;
    din_valid_1_28 <= out_new_pkt | hash_out_valid_filter_1_28;
    din_valid_1_28_r1 <= din_valid_1_28;
    din_valid_1_28_r2 <= din_valid_1_28_r1;

    din_1_28.data <= hash_out_valid_filter_1_28 ? hash_out_1_28 : 0;
    din_1_28.last <= out_new_pkt;
    din_1_28.bucket <= 1;


    din_1_28_r1 <= din_1_28;
    din_1_28_r2 <= din_1_28_r1;
    din_valid_1_29 <= out_new_pkt | hash_out_valid_filter_1_29;
    din_valid_1_29_r1 <= din_valid_1_29;
    din_valid_1_29_r2 <= din_valid_1_29_r1;

    din_1_29.data <= hash_out_valid_filter_1_29 ? hash_out_1_29 : 0;
    din_1_29.last <= out_new_pkt;
    din_1_29.bucket <= 1;


    din_1_29_r1 <= din_1_29;
    din_1_29_r2 <= din_1_29_r1;
    din_valid_1_30 <= out_new_pkt | hash_out_valid_filter_1_30;
    din_valid_1_30_r1 <= din_valid_1_30;
    din_valid_1_30_r2 <= din_valid_1_30_r1;

    din_1_30.data <= hash_out_valid_filter_1_30 ? hash_out_1_30 : 0;
    din_1_30.last <= out_new_pkt;
    din_1_30.bucket <= 1;


    din_1_30_r1 <= din_1_30;
    din_1_30_r2 <= din_1_30_r1;
    din_valid_1_31 <= out_new_pkt | hash_out_valid_filter_1_31;
    din_valid_1_31_r1 <= din_valid_1_31;
    din_valid_1_31_r2 <= din_valid_1_31_r1;

    din_1_31.data <= hash_out_valid_filter_1_31 ? hash_out_1_31 : 0;
    din_1_31.last <= out_new_pkt;
    din_1_31.bucket <= 1;


    din_1_31_r1 <= din_1_31;
    din_1_31_r2 <= din_1_31_r1;
    din_valid_2_0 <= out_new_pkt | hash_out_valid_filter_2_0;
    din_valid_2_0_r1 <= din_valid_2_0;
    din_valid_2_0_r2 <= din_valid_2_0_r1;

    din_2_0.data <= hash_out_valid_filter_2_0 ? hash_out_2_0 : 0;
    din_2_0.last <= out_new_pkt;
    din_2_0.bucket <= 2;


    din_2_0_r1 <= din_2_0;
    din_2_0_r2 <= din_2_0_r1;
    din_valid_2_1 <= out_new_pkt | hash_out_valid_filter_2_1;
    din_valid_2_1_r1 <= din_valid_2_1;
    din_valid_2_1_r2 <= din_valid_2_1_r1;

    din_2_1.data <= hash_out_valid_filter_2_1 ? hash_out_2_1 : 0;
    din_2_1.last <= out_new_pkt;
    din_2_1.bucket <= 2;


    din_2_1_r1 <= din_2_1;
    din_2_1_r2 <= din_2_1_r1;
    din_valid_2_2 <= out_new_pkt | hash_out_valid_filter_2_2;
    din_valid_2_2_r1 <= din_valid_2_2;
    din_valid_2_2_r2 <= din_valid_2_2_r1;

    din_2_2.data <= hash_out_valid_filter_2_2 ? hash_out_2_2 : 0;
    din_2_2.last <= out_new_pkt;
    din_2_2.bucket <= 2;


    din_2_2_r1 <= din_2_2;
    din_2_2_r2 <= din_2_2_r1;
    din_valid_2_3 <= out_new_pkt | hash_out_valid_filter_2_3;
    din_valid_2_3_r1 <= din_valid_2_3;
    din_valid_2_3_r2 <= din_valid_2_3_r1;

    din_2_3.data <= hash_out_valid_filter_2_3 ? hash_out_2_3 : 0;
    din_2_3.last <= out_new_pkt;
    din_2_3.bucket <= 2;


    din_2_3_r1 <= din_2_3;
    din_2_3_r2 <= din_2_3_r1;
    din_valid_2_4 <= out_new_pkt | hash_out_valid_filter_2_4;
    din_valid_2_4_r1 <= din_valid_2_4;
    din_valid_2_4_r2 <= din_valid_2_4_r1;

    din_2_4.data <= hash_out_valid_filter_2_4 ? hash_out_2_4 : 0;
    din_2_4.last <= out_new_pkt;
    din_2_4.bucket <= 2;


    din_2_4_r1 <= din_2_4;
    din_2_4_r2 <= din_2_4_r1;
    din_valid_2_5 <= out_new_pkt | hash_out_valid_filter_2_5;
    din_valid_2_5_r1 <= din_valid_2_5;
    din_valid_2_5_r2 <= din_valid_2_5_r1;

    din_2_5.data <= hash_out_valid_filter_2_5 ? hash_out_2_5 : 0;
    din_2_5.last <= out_new_pkt;
    din_2_5.bucket <= 2;


    din_2_5_r1 <= din_2_5;
    din_2_5_r2 <= din_2_5_r1;
    din_valid_2_6 <= out_new_pkt | hash_out_valid_filter_2_6;
    din_valid_2_6_r1 <= din_valid_2_6;
    din_valid_2_6_r2 <= din_valid_2_6_r1;

    din_2_6.data <= hash_out_valid_filter_2_6 ? hash_out_2_6 : 0;
    din_2_6.last <= out_new_pkt;
    din_2_6.bucket <= 2;


    din_2_6_r1 <= din_2_6;
    din_2_6_r2 <= din_2_6_r1;
    din_valid_2_7 <= out_new_pkt | hash_out_valid_filter_2_7;
    din_valid_2_7_r1 <= din_valid_2_7;
    din_valid_2_7_r2 <= din_valid_2_7_r1;

    din_2_7.data <= hash_out_valid_filter_2_7 ? hash_out_2_7 : 0;
    din_2_7.last <= out_new_pkt;
    din_2_7.bucket <= 2;


    din_2_7_r1 <= din_2_7;
    din_2_7_r2 <= din_2_7_r1;
    din_valid_2_8 <= out_new_pkt | hash_out_valid_filter_2_8;
    din_valid_2_8_r1 <= din_valid_2_8;
    din_valid_2_8_r2 <= din_valid_2_8_r1;

    din_2_8.data <= hash_out_valid_filter_2_8 ? hash_out_2_8 : 0;
    din_2_8.last <= out_new_pkt;
    din_2_8.bucket <= 2;


    din_2_8_r1 <= din_2_8;
    din_2_8_r2 <= din_2_8_r1;
    din_valid_2_9 <= out_new_pkt | hash_out_valid_filter_2_9;
    din_valid_2_9_r1 <= din_valid_2_9;
    din_valid_2_9_r2 <= din_valid_2_9_r1;

    din_2_9.data <= hash_out_valid_filter_2_9 ? hash_out_2_9 : 0;
    din_2_9.last <= out_new_pkt;
    din_2_9.bucket <= 2;


    din_2_9_r1 <= din_2_9;
    din_2_9_r2 <= din_2_9_r1;
    din_valid_2_10 <= out_new_pkt | hash_out_valid_filter_2_10;
    din_valid_2_10_r1 <= din_valid_2_10;
    din_valid_2_10_r2 <= din_valid_2_10_r1;

    din_2_10.data <= hash_out_valid_filter_2_10 ? hash_out_2_10 : 0;
    din_2_10.last <= out_new_pkt;
    din_2_10.bucket <= 2;


    din_2_10_r1 <= din_2_10;
    din_2_10_r2 <= din_2_10_r1;
    din_valid_2_11 <= out_new_pkt | hash_out_valid_filter_2_11;
    din_valid_2_11_r1 <= din_valid_2_11;
    din_valid_2_11_r2 <= din_valid_2_11_r1;

    din_2_11.data <= hash_out_valid_filter_2_11 ? hash_out_2_11 : 0;
    din_2_11.last <= out_new_pkt;
    din_2_11.bucket <= 2;


    din_2_11_r1 <= din_2_11;
    din_2_11_r2 <= din_2_11_r1;
    din_valid_2_12 <= out_new_pkt | hash_out_valid_filter_2_12;
    din_valid_2_12_r1 <= din_valid_2_12;
    din_valid_2_12_r2 <= din_valid_2_12_r1;

    din_2_12.data <= hash_out_valid_filter_2_12 ? hash_out_2_12 : 0;
    din_2_12.last <= out_new_pkt;
    din_2_12.bucket <= 2;


    din_2_12_r1 <= din_2_12;
    din_2_12_r2 <= din_2_12_r1;
    din_valid_2_13 <= out_new_pkt | hash_out_valid_filter_2_13;
    din_valid_2_13_r1 <= din_valid_2_13;
    din_valid_2_13_r2 <= din_valid_2_13_r1;

    din_2_13.data <= hash_out_valid_filter_2_13 ? hash_out_2_13 : 0;
    din_2_13.last <= out_new_pkt;
    din_2_13.bucket <= 2;


    din_2_13_r1 <= din_2_13;
    din_2_13_r2 <= din_2_13_r1;
    din_valid_2_14 <= out_new_pkt | hash_out_valid_filter_2_14;
    din_valid_2_14_r1 <= din_valid_2_14;
    din_valid_2_14_r2 <= din_valid_2_14_r1;

    din_2_14.data <= hash_out_valid_filter_2_14 ? hash_out_2_14 : 0;
    din_2_14.last <= out_new_pkt;
    din_2_14.bucket <= 2;


    din_2_14_r1 <= din_2_14;
    din_2_14_r2 <= din_2_14_r1;
    din_valid_2_15 <= out_new_pkt | hash_out_valid_filter_2_15;
    din_valid_2_15_r1 <= din_valid_2_15;
    din_valid_2_15_r2 <= din_valid_2_15_r1;

    din_2_15.data <= hash_out_valid_filter_2_15 ? hash_out_2_15 : 0;
    din_2_15.last <= out_new_pkt;
    din_2_15.bucket <= 2;


    din_2_15_r1 <= din_2_15;
    din_2_15_r2 <= din_2_15_r1;
    din_valid_2_16 <= out_new_pkt | hash_out_valid_filter_2_16;
    din_valid_2_16_r1 <= din_valid_2_16;
    din_valid_2_16_r2 <= din_valid_2_16_r1;

    din_2_16.data <= hash_out_valid_filter_2_16 ? hash_out_2_16 : 0;
    din_2_16.last <= out_new_pkt;
    din_2_16.bucket <= 2;


    din_2_16_r1 <= din_2_16;
    din_2_16_r2 <= din_2_16_r1;
    din_valid_2_17 <= out_new_pkt | hash_out_valid_filter_2_17;
    din_valid_2_17_r1 <= din_valid_2_17;
    din_valid_2_17_r2 <= din_valid_2_17_r1;

    din_2_17.data <= hash_out_valid_filter_2_17 ? hash_out_2_17 : 0;
    din_2_17.last <= out_new_pkt;
    din_2_17.bucket <= 2;


    din_2_17_r1 <= din_2_17;
    din_2_17_r2 <= din_2_17_r1;
    din_valid_2_18 <= out_new_pkt | hash_out_valid_filter_2_18;
    din_valid_2_18_r1 <= din_valid_2_18;
    din_valid_2_18_r2 <= din_valid_2_18_r1;

    din_2_18.data <= hash_out_valid_filter_2_18 ? hash_out_2_18 : 0;
    din_2_18.last <= out_new_pkt;
    din_2_18.bucket <= 2;


    din_2_18_r1 <= din_2_18;
    din_2_18_r2 <= din_2_18_r1;
    din_valid_2_19 <= out_new_pkt | hash_out_valid_filter_2_19;
    din_valid_2_19_r1 <= din_valid_2_19;
    din_valid_2_19_r2 <= din_valid_2_19_r1;

    din_2_19.data <= hash_out_valid_filter_2_19 ? hash_out_2_19 : 0;
    din_2_19.last <= out_new_pkt;
    din_2_19.bucket <= 2;


    din_2_19_r1 <= din_2_19;
    din_2_19_r2 <= din_2_19_r1;
    din_valid_2_20 <= out_new_pkt | hash_out_valid_filter_2_20;
    din_valid_2_20_r1 <= din_valid_2_20;
    din_valid_2_20_r2 <= din_valid_2_20_r1;

    din_2_20.data <= hash_out_valid_filter_2_20 ? hash_out_2_20 : 0;
    din_2_20.last <= out_new_pkt;
    din_2_20.bucket <= 2;


    din_2_20_r1 <= din_2_20;
    din_2_20_r2 <= din_2_20_r1;
    din_valid_2_21 <= out_new_pkt | hash_out_valid_filter_2_21;
    din_valid_2_21_r1 <= din_valid_2_21;
    din_valid_2_21_r2 <= din_valid_2_21_r1;

    din_2_21.data <= hash_out_valid_filter_2_21 ? hash_out_2_21 : 0;
    din_2_21.last <= out_new_pkt;
    din_2_21.bucket <= 2;


    din_2_21_r1 <= din_2_21;
    din_2_21_r2 <= din_2_21_r1;
    din_valid_2_22 <= out_new_pkt | hash_out_valid_filter_2_22;
    din_valid_2_22_r1 <= din_valid_2_22;
    din_valid_2_22_r2 <= din_valid_2_22_r1;

    din_2_22.data <= hash_out_valid_filter_2_22 ? hash_out_2_22 : 0;
    din_2_22.last <= out_new_pkt;
    din_2_22.bucket <= 2;


    din_2_22_r1 <= din_2_22;
    din_2_22_r2 <= din_2_22_r1;
    din_valid_2_23 <= out_new_pkt | hash_out_valid_filter_2_23;
    din_valid_2_23_r1 <= din_valid_2_23;
    din_valid_2_23_r2 <= din_valid_2_23_r1;

    din_2_23.data <= hash_out_valid_filter_2_23 ? hash_out_2_23 : 0;
    din_2_23.last <= out_new_pkt;
    din_2_23.bucket <= 2;


    din_2_23_r1 <= din_2_23;
    din_2_23_r2 <= din_2_23_r1;
    din_valid_2_24 <= out_new_pkt | hash_out_valid_filter_2_24;
    din_valid_2_24_r1 <= din_valid_2_24;
    din_valid_2_24_r2 <= din_valid_2_24_r1;

    din_2_24.data <= hash_out_valid_filter_2_24 ? hash_out_2_24 : 0;
    din_2_24.last <= out_new_pkt;
    din_2_24.bucket <= 2;


    din_2_24_r1 <= din_2_24;
    din_2_24_r2 <= din_2_24_r1;
    din_valid_2_25 <= out_new_pkt | hash_out_valid_filter_2_25;
    din_valid_2_25_r1 <= din_valid_2_25;
    din_valid_2_25_r2 <= din_valid_2_25_r1;

    din_2_25.data <= hash_out_valid_filter_2_25 ? hash_out_2_25 : 0;
    din_2_25.last <= out_new_pkt;
    din_2_25.bucket <= 2;


    din_2_25_r1 <= din_2_25;
    din_2_25_r2 <= din_2_25_r1;
    din_valid_2_26 <= out_new_pkt | hash_out_valid_filter_2_26;
    din_valid_2_26_r1 <= din_valid_2_26;
    din_valid_2_26_r2 <= din_valid_2_26_r1;

    din_2_26.data <= hash_out_valid_filter_2_26 ? hash_out_2_26 : 0;
    din_2_26.last <= out_new_pkt;
    din_2_26.bucket <= 2;


    din_2_26_r1 <= din_2_26;
    din_2_26_r2 <= din_2_26_r1;
    din_valid_2_27 <= out_new_pkt | hash_out_valid_filter_2_27;
    din_valid_2_27_r1 <= din_valid_2_27;
    din_valid_2_27_r2 <= din_valid_2_27_r1;

    din_2_27.data <= hash_out_valid_filter_2_27 ? hash_out_2_27 : 0;
    din_2_27.last <= out_new_pkt;
    din_2_27.bucket <= 2;


    din_2_27_r1 <= din_2_27;
    din_2_27_r2 <= din_2_27_r1;
    din_valid_2_28 <= out_new_pkt | hash_out_valid_filter_2_28;
    din_valid_2_28_r1 <= din_valid_2_28;
    din_valid_2_28_r2 <= din_valid_2_28_r1;

    din_2_28.data <= hash_out_valid_filter_2_28 ? hash_out_2_28 : 0;
    din_2_28.last <= out_new_pkt;
    din_2_28.bucket <= 2;


    din_2_28_r1 <= din_2_28;
    din_2_28_r2 <= din_2_28_r1;
    din_valid_2_29 <= out_new_pkt | hash_out_valid_filter_2_29;
    din_valid_2_29_r1 <= din_valid_2_29;
    din_valid_2_29_r2 <= din_valid_2_29_r1;

    din_2_29.data <= hash_out_valid_filter_2_29 ? hash_out_2_29 : 0;
    din_2_29.last <= out_new_pkt;
    din_2_29.bucket <= 2;


    din_2_29_r1 <= din_2_29;
    din_2_29_r2 <= din_2_29_r1;
    din_valid_2_30 <= out_new_pkt | hash_out_valid_filter_2_30;
    din_valid_2_30_r1 <= din_valid_2_30;
    din_valid_2_30_r2 <= din_valid_2_30_r1;

    din_2_30.data <= hash_out_valid_filter_2_30 ? hash_out_2_30 : 0;
    din_2_30.last <= out_new_pkt;
    din_2_30.bucket <= 2;


    din_2_30_r1 <= din_2_30;
    din_2_30_r2 <= din_2_30_r1;
    din_valid_2_31 <= out_new_pkt | hash_out_valid_filter_2_31;
    din_valid_2_31_r1 <= din_valid_2_31;
    din_valid_2_31_r2 <= din_valid_2_31_r1;

    din_2_31.data <= hash_out_valid_filter_2_31 ? hash_out_2_31 : 0;
    din_2_31.last <= out_new_pkt;
    din_2_31.bucket <= 2;


    din_2_31_r1 <= din_2_31;
    din_2_31_r2 <= din_2_31_r1;
    din_valid_3_0 <= out_new_pkt | hash_out_valid_filter_3_0;
    din_valid_3_0_r1 <= din_valid_3_0;
    din_valid_3_0_r2 <= din_valid_3_0_r1;

    din_3_0.data <= hash_out_valid_filter_3_0 ? hash_out_3_0 : 0;
    din_3_0.last <= out_new_pkt;
    din_3_0.bucket <= 3;


    din_3_0_r1 <= din_3_0;
    din_3_0_r2 <= din_3_0_r1;
    din_valid_3_1 <= out_new_pkt | hash_out_valid_filter_3_1;
    din_valid_3_1_r1 <= din_valid_3_1;
    din_valid_3_1_r2 <= din_valid_3_1_r1;

    din_3_1.data <= hash_out_valid_filter_3_1 ? hash_out_3_1 : 0;
    din_3_1.last <= out_new_pkt;
    din_3_1.bucket <= 3;


    din_3_1_r1 <= din_3_1;
    din_3_1_r2 <= din_3_1_r1;
    din_valid_3_2 <= out_new_pkt | hash_out_valid_filter_3_2;
    din_valid_3_2_r1 <= din_valid_3_2;
    din_valid_3_2_r2 <= din_valid_3_2_r1;

    din_3_2.data <= hash_out_valid_filter_3_2 ? hash_out_3_2 : 0;
    din_3_2.last <= out_new_pkt;
    din_3_2.bucket <= 3;


    din_3_2_r1 <= din_3_2;
    din_3_2_r2 <= din_3_2_r1;
    din_valid_3_3 <= out_new_pkt | hash_out_valid_filter_3_3;
    din_valid_3_3_r1 <= din_valid_3_3;
    din_valid_3_3_r2 <= din_valid_3_3_r1;

    din_3_3.data <= hash_out_valid_filter_3_3 ? hash_out_3_3 : 0;
    din_3_3.last <= out_new_pkt;
    din_3_3.bucket <= 3;


    din_3_3_r1 <= din_3_3;
    din_3_3_r2 <= din_3_3_r1;
    din_valid_3_4 <= out_new_pkt | hash_out_valid_filter_3_4;
    din_valid_3_4_r1 <= din_valid_3_4;
    din_valid_3_4_r2 <= din_valid_3_4_r1;

    din_3_4.data <= hash_out_valid_filter_3_4 ? hash_out_3_4 : 0;
    din_3_4.last <= out_new_pkt;
    din_3_4.bucket <= 3;


    din_3_4_r1 <= din_3_4;
    din_3_4_r2 <= din_3_4_r1;
    din_valid_3_5 <= out_new_pkt | hash_out_valid_filter_3_5;
    din_valid_3_5_r1 <= din_valid_3_5;
    din_valid_3_5_r2 <= din_valid_3_5_r1;

    din_3_5.data <= hash_out_valid_filter_3_5 ? hash_out_3_5 : 0;
    din_3_5.last <= out_new_pkt;
    din_3_5.bucket <= 3;


    din_3_5_r1 <= din_3_5;
    din_3_5_r2 <= din_3_5_r1;
    din_valid_3_6 <= out_new_pkt | hash_out_valid_filter_3_6;
    din_valid_3_6_r1 <= din_valid_3_6;
    din_valid_3_6_r2 <= din_valid_3_6_r1;

    din_3_6.data <= hash_out_valid_filter_3_6 ? hash_out_3_6 : 0;
    din_3_6.last <= out_new_pkt;
    din_3_6.bucket <= 3;


    din_3_6_r1 <= din_3_6;
    din_3_6_r2 <= din_3_6_r1;
    din_valid_3_7 <= out_new_pkt | hash_out_valid_filter_3_7;
    din_valid_3_7_r1 <= din_valid_3_7;
    din_valid_3_7_r2 <= din_valid_3_7_r1;

    din_3_7.data <= hash_out_valid_filter_3_7 ? hash_out_3_7 : 0;
    din_3_7.last <= out_new_pkt;
    din_3_7.bucket <= 3;


    din_3_7_r1 <= din_3_7;
    din_3_7_r2 <= din_3_7_r1;
    din_valid_3_8 <= out_new_pkt | hash_out_valid_filter_3_8;
    din_valid_3_8_r1 <= din_valid_3_8;
    din_valid_3_8_r2 <= din_valid_3_8_r1;

    din_3_8.data <= hash_out_valid_filter_3_8 ? hash_out_3_8 : 0;
    din_3_8.last <= out_new_pkt;
    din_3_8.bucket <= 3;


    din_3_8_r1 <= din_3_8;
    din_3_8_r2 <= din_3_8_r1;
    din_valid_3_9 <= out_new_pkt | hash_out_valid_filter_3_9;
    din_valid_3_9_r1 <= din_valid_3_9;
    din_valid_3_9_r2 <= din_valid_3_9_r1;

    din_3_9.data <= hash_out_valid_filter_3_9 ? hash_out_3_9 : 0;
    din_3_9.last <= out_new_pkt;
    din_3_9.bucket <= 3;


    din_3_9_r1 <= din_3_9;
    din_3_9_r2 <= din_3_9_r1;
    din_valid_3_10 <= out_new_pkt | hash_out_valid_filter_3_10;
    din_valid_3_10_r1 <= din_valid_3_10;
    din_valid_3_10_r2 <= din_valid_3_10_r1;

    din_3_10.data <= hash_out_valid_filter_3_10 ? hash_out_3_10 : 0;
    din_3_10.last <= out_new_pkt;
    din_3_10.bucket <= 3;


    din_3_10_r1 <= din_3_10;
    din_3_10_r2 <= din_3_10_r1;
    din_valid_3_11 <= out_new_pkt | hash_out_valid_filter_3_11;
    din_valid_3_11_r1 <= din_valid_3_11;
    din_valid_3_11_r2 <= din_valid_3_11_r1;

    din_3_11.data <= hash_out_valid_filter_3_11 ? hash_out_3_11 : 0;
    din_3_11.last <= out_new_pkt;
    din_3_11.bucket <= 3;


    din_3_11_r1 <= din_3_11;
    din_3_11_r2 <= din_3_11_r1;
    din_valid_3_12 <= out_new_pkt | hash_out_valid_filter_3_12;
    din_valid_3_12_r1 <= din_valid_3_12;
    din_valid_3_12_r2 <= din_valid_3_12_r1;

    din_3_12.data <= hash_out_valid_filter_3_12 ? hash_out_3_12 : 0;
    din_3_12.last <= out_new_pkt;
    din_3_12.bucket <= 3;


    din_3_12_r1 <= din_3_12;
    din_3_12_r2 <= din_3_12_r1;
    din_valid_3_13 <= out_new_pkt | hash_out_valid_filter_3_13;
    din_valid_3_13_r1 <= din_valid_3_13;
    din_valid_3_13_r2 <= din_valid_3_13_r1;

    din_3_13.data <= hash_out_valid_filter_3_13 ? hash_out_3_13 : 0;
    din_3_13.last <= out_new_pkt;
    din_3_13.bucket <= 3;


    din_3_13_r1 <= din_3_13;
    din_3_13_r2 <= din_3_13_r1;
    din_valid_3_14 <= out_new_pkt | hash_out_valid_filter_3_14;
    din_valid_3_14_r1 <= din_valid_3_14;
    din_valid_3_14_r2 <= din_valid_3_14_r1;

    din_3_14.data <= hash_out_valid_filter_3_14 ? hash_out_3_14 : 0;
    din_3_14.last <= out_new_pkt;
    din_3_14.bucket <= 3;


    din_3_14_r1 <= din_3_14;
    din_3_14_r2 <= din_3_14_r1;
    din_valid_3_15 <= out_new_pkt | hash_out_valid_filter_3_15;
    din_valid_3_15_r1 <= din_valid_3_15;
    din_valid_3_15_r2 <= din_valid_3_15_r1;

    din_3_15.data <= hash_out_valid_filter_3_15 ? hash_out_3_15 : 0;
    din_3_15.last <= out_new_pkt;
    din_3_15.bucket <= 3;


    din_3_15_r1 <= din_3_15;
    din_3_15_r2 <= din_3_15_r1;
    din_valid_3_16 <= out_new_pkt | hash_out_valid_filter_3_16;
    din_valid_3_16_r1 <= din_valid_3_16;
    din_valid_3_16_r2 <= din_valid_3_16_r1;

    din_3_16.data <= hash_out_valid_filter_3_16 ? hash_out_3_16 : 0;
    din_3_16.last <= out_new_pkt;
    din_3_16.bucket <= 3;


    din_3_16_r1 <= din_3_16;
    din_3_16_r2 <= din_3_16_r1;
    din_valid_3_17 <= out_new_pkt | hash_out_valid_filter_3_17;
    din_valid_3_17_r1 <= din_valid_3_17;
    din_valid_3_17_r2 <= din_valid_3_17_r1;

    din_3_17.data <= hash_out_valid_filter_3_17 ? hash_out_3_17 : 0;
    din_3_17.last <= out_new_pkt;
    din_3_17.bucket <= 3;


    din_3_17_r1 <= din_3_17;
    din_3_17_r2 <= din_3_17_r1;
    din_valid_3_18 <= out_new_pkt | hash_out_valid_filter_3_18;
    din_valid_3_18_r1 <= din_valid_3_18;
    din_valid_3_18_r2 <= din_valid_3_18_r1;

    din_3_18.data <= hash_out_valid_filter_3_18 ? hash_out_3_18 : 0;
    din_3_18.last <= out_new_pkt;
    din_3_18.bucket <= 3;


    din_3_18_r1 <= din_3_18;
    din_3_18_r2 <= din_3_18_r1;
    din_valid_3_19 <= out_new_pkt | hash_out_valid_filter_3_19;
    din_valid_3_19_r1 <= din_valid_3_19;
    din_valid_3_19_r2 <= din_valid_3_19_r1;

    din_3_19.data <= hash_out_valid_filter_3_19 ? hash_out_3_19 : 0;
    din_3_19.last <= out_new_pkt;
    din_3_19.bucket <= 3;


    din_3_19_r1 <= din_3_19;
    din_3_19_r2 <= din_3_19_r1;
    din_valid_3_20 <= out_new_pkt | hash_out_valid_filter_3_20;
    din_valid_3_20_r1 <= din_valid_3_20;
    din_valid_3_20_r2 <= din_valid_3_20_r1;

    din_3_20.data <= hash_out_valid_filter_3_20 ? hash_out_3_20 : 0;
    din_3_20.last <= out_new_pkt;
    din_3_20.bucket <= 3;


    din_3_20_r1 <= din_3_20;
    din_3_20_r2 <= din_3_20_r1;
    din_valid_3_21 <= out_new_pkt | hash_out_valid_filter_3_21;
    din_valid_3_21_r1 <= din_valid_3_21;
    din_valid_3_21_r2 <= din_valid_3_21_r1;

    din_3_21.data <= hash_out_valid_filter_3_21 ? hash_out_3_21 : 0;
    din_3_21.last <= out_new_pkt;
    din_3_21.bucket <= 3;


    din_3_21_r1 <= din_3_21;
    din_3_21_r2 <= din_3_21_r1;
    din_valid_3_22 <= out_new_pkt | hash_out_valid_filter_3_22;
    din_valid_3_22_r1 <= din_valid_3_22;
    din_valid_3_22_r2 <= din_valid_3_22_r1;

    din_3_22.data <= hash_out_valid_filter_3_22 ? hash_out_3_22 : 0;
    din_3_22.last <= out_new_pkt;
    din_3_22.bucket <= 3;


    din_3_22_r1 <= din_3_22;
    din_3_22_r2 <= din_3_22_r1;
    din_valid_3_23 <= out_new_pkt | hash_out_valid_filter_3_23;
    din_valid_3_23_r1 <= din_valid_3_23;
    din_valid_3_23_r2 <= din_valid_3_23_r1;

    din_3_23.data <= hash_out_valid_filter_3_23 ? hash_out_3_23 : 0;
    din_3_23.last <= out_new_pkt;
    din_3_23.bucket <= 3;


    din_3_23_r1 <= din_3_23;
    din_3_23_r2 <= din_3_23_r1;
    din_valid_3_24 <= out_new_pkt | hash_out_valid_filter_3_24;
    din_valid_3_24_r1 <= din_valid_3_24;
    din_valid_3_24_r2 <= din_valid_3_24_r1;

    din_3_24.data <= hash_out_valid_filter_3_24 ? hash_out_3_24 : 0;
    din_3_24.last <= out_new_pkt;
    din_3_24.bucket <= 3;


    din_3_24_r1 <= din_3_24;
    din_3_24_r2 <= din_3_24_r1;
    din_valid_3_25 <= out_new_pkt | hash_out_valid_filter_3_25;
    din_valid_3_25_r1 <= din_valid_3_25;
    din_valid_3_25_r2 <= din_valid_3_25_r1;

    din_3_25.data <= hash_out_valid_filter_3_25 ? hash_out_3_25 : 0;
    din_3_25.last <= out_new_pkt;
    din_3_25.bucket <= 3;


    din_3_25_r1 <= din_3_25;
    din_3_25_r2 <= din_3_25_r1;
    din_valid_3_26 <= out_new_pkt | hash_out_valid_filter_3_26;
    din_valid_3_26_r1 <= din_valid_3_26;
    din_valid_3_26_r2 <= din_valid_3_26_r1;

    din_3_26.data <= hash_out_valid_filter_3_26 ? hash_out_3_26 : 0;
    din_3_26.last <= out_new_pkt;
    din_3_26.bucket <= 3;


    din_3_26_r1 <= din_3_26;
    din_3_26_r2 <= din_3_26_r1;
    din_valid_3_27 <= out_new_pkt | hash_out_valid_filter_3_27;
    din_valid_3_27_r1 <= din_valid_3_27;
    din_valid_3_27_r2 <= din_valid_3_27_r1;

    din_3_27.data <= hash_out_valid_filter_3_27 ? hash_out_3_27 : 0;
    din_3_27.last <= out_new_pkt;
    din_3_27.bucket <= 3;


    din_3_27_r1 <= din_3_27;
    din_3_27_r2 <= din_3_27_r1;
    din_valid_3_28 <= out_new_pkt | hash_out_valid_filter_3_28;
    din_valid_3_28_r1 <= din_valid_3_28;
    din_valid_3_28_r2 <= din_valid_3_28_r1;

    din_3_28.data <= hash_out_valid_filter_3_28 ? hash_out_3_28 : 0;
    din_3_28.last <= out_new_pkt;
    din_3_28.bucket <= 3;


    din_3_28_r1 <= din_3_28;
    din_3_28_r2 <= din_3_28_r1;
    din_valid_3_29 <= out_new_pkt | hash_out_valid_filter_3_29;
    din_valid_3_29_r1 <= din_valid_3_29;
    din_valid_3_29_r2 <= din_valid_3_29_r1;

    din_3_29.data <= hash_out_valid_filter_3_29 ? hash_out_3_29 : 0;
    din_3_29.last <= out_new_pkt;
    din_3_29.bucket <= 3;


    din_3_29_r1 <= din_3_29;
    din_3_29_r2 <= din_3_29_r1;
    din_valid_3_30 <= out_new_pkt | hash_out_valid_filter_3_30;
    din_valid_3_30_r1 <= din_valid_3_30;
    din_valid_3_30_r2 <= din_valid_3_30_r1;

    din_3_30.data <= hash_out_valid_filter_3_30 ? hash_out_3_30 : 0;
    din_3_30.last <= out_new_pkt;
    din_3_30.bucket <= 3;


    din_3_30_r1 <= din_3_30;
    din_3_30_r2 <= din_3_30_r1;
    din_valid_3_31 <= out_new_pkt | hash_out_valid_filter_3_31;
    din_valid_3_31_r1 <= din_valid_3_31;
    din_valid_3_31_r2 <= din_valid_3_31_r1;

    din_3_31.data <= hash_out_valid_filter_3_31 ? hash_out_3_31 : 0;
    din_3_31.last <= out_new_pkt;
    din_3_31.bucket <= 3;


    din_3_31_r1 <= din_3_31;
    din_3_31_r2 <= din_3_31_r1;
    din_valid_4_0 <= out_new_pkt | hash_out_valid_filter_4_0;
    din_valid_4_0_r1 <= din_valid_4_0;
    din_valid_4_0_r2 <= din_valid_4_0_r1;

    din_4_0.data <= hash_out_valid_filter_4_0 ? hash_out_4_0 : 0;
    din_4_0.last <= out_new_pkt;
    din_4_0.bucket <= 4;


    din_4_0_r1 <= din_4_0;
    din_4_0_r2 <= din_4_0_r1;
    din_valid_4_1 <= out_new_pkt | hash_out_valid_filter_4_1;
    din_valid_4_1_r1 <= din_valid_4_1;
    din_valid_4_1_r2 <= din_valid_4_1_r1;

    din_4_1.data <= hash_out_valid_filter_4_1 ? hash_out_4_1 : 0;
    din_4_1.last <= out_new_pkt;
    din_4_1.bucket <= 4;


    din_4_1_r1 <= din_4_1;
    din_4_1_r2 <= din_4_1_r1;
    din_valid_4_2 <= out_new_pkt | hash_out_valid_filter_4_2;
    din_valid_4_2_r1 <= din_valid_4_2;
    din_valid_4_2_r2 <= din_valid_4_2_r1;

    din_4_2.data <= hash_out_valid_filter_4_2 ? hash_out_4_2 : 0;
    din_4_2.last <= out_new_pkt;
    din_4_2.bucket <= 4;


    din_4_2_r1 <= din_4_2;
    din_4_2_r2 <= din_4_2_r1;
    din_valid_4_3 <= out_new_pkt | hash_out_valid_filter_4_3;
    din_valid_4_3_r1 <= din_valid_4_3;
    din_valid_4_3_r2 <= din_valid_4_3_r1;

    din_4_3.data <= hash_out_valid_filter_4_3 ? hash_out_4_3 : 0;
    din_4_3.last <= out_new_pkt;
    din_4_3.bucket <= 4;


    din_4_3_r1 <= din_4_3;
    din_4_3_r2 <= din_4_3_r1;
    din_valid_4_4 <= out_new_pkt | hash_out_valid_filter_4_4;
    din_valid_4_4_r1 <= din_valid_4_4;
    din_valid_4_4_r2 <= din_valid_4_4_r1;

    din_4_4.data <= hash_out_valid_filter_4_4 ? hash_out_4_4 : 0;
    din_4_4.last <= out_new_pkt;
    din_4_4.bucket <= 4;


    din_4_4_r1 <= din_4_4;
    din_4_4_r2 <= din_4_4_r1;
    din_valid_4_5 <= out_new_pkt | hash_out_valid_filter_4_5;
    din_valid_4_5_r1 <= din_valid_4_5;
    din_valid_4_5_r2 <= din_valid_4_5_r1;

    din_4_5.data <= hash_out_valid_filter_4_5 ? hash_out_4_5 : 0;
    din_4_5.last <= out_new_pkt;
    din_4_5.bucket <= 4;


    din_4_5_r1 <= din_4_5;
    din_4_5_r2 <= din_4_5_r1;
    din_valid_4_6 <= out_new_pkt | hash_out_valid_filter_4_6;
    din_valid_4_6_r1 <= din_valid_4_6;
    din_valid_4_6_r2 <= din_valid_4_6_r1;

    din_4_6.data <= hash_out_valid_filter_4_6 ? hash_out_4_6 : 0;
    din_4_6.last <= out_new_pkt;
    din_4_6.bucket <= 4;


    din_4_6_r1 <= din_4_6;
    din_4_6_r2 <= din_4_6_r1;
    din_valid_4_7 <= out_new_pkt | hash_out_valid_filter_4_7;
    din_valid_4_7_r1 <= din_valid_4_7;
    din_valid_4_7_r2 <= din_valid_4_7_r1;

    din_4_7.data <= hash_out_valid_filter_4_7 ? hash_out_4_7 : 0;
    din_4_7.last <= out_new_pkt;
    din_4_7.bucket <= 4;


    din_4_7_r1 <= din_4_7;
    din_4_7_r2 <= din_4_7_r1;
    din_valid_4_8 <= out_new_pkt | hash_out_valid_filter_4_8;
    din_valid_4_8_r1 <= din_valid_4_8;
    din_valid_4_8_r2 <= din_valid_4_8_r1;

    din_4_8.data <= hash_out_valid_filter_4_8 ? hash_out_4_8 : 0;
    din_4_8.last <= out_new_pkt;
    din_4_8.bucket <= 4;


    din_4_8_r1 <= din_4_8;
    din_4_8_r2 <= din_4_8_r1;
    din_valid_4_9 <= out_new_pkt | hash_out_valid_filter_4_9;
    din_valid_4_9_r1 <= din_valid_4_9;
    din_valid_4_9_r2 <= din_valid_4_9_r1;

    din_4_9.data <= hash_out_valid_filter_4_9 ? hash_out_4_9 : 0;
    din_4_9.last <= out_new_pkt;
    din_4_9.bucket <= 4;


    din_4_9_r1 <= din_4_9;
    din_4_9_r2 <= din_4_9_r1;
    din_valid_4_10 <= out_new_pkt | hash_out_valid_filter_4_10;
    din_valid_4_10_r1 <= din_valid_4_10;
    din_valid_4_10_r2 <= din_valid_4_10_r1;

    din_4_10.data <= hash_out_valid_filter_4_10 ? hash_out_4_10 : 0;
    din_4_10.last <= out_new_pkt;
    din_4_10.bucket <= 4;


    din_4_10_r1 <= din_4_10;
    din_4_10_r2 <= din_4_10_r1;
    din_valid_4_11 <= out_new_pkt | hash_out_valid_filter_4_11;
    din_valid_4_11_r1 <= din_valid_4_11;
    din_valid_4_11_r2 <= din_valid_4_11_r1;

    din_4_11.data <= hash_out_valid_filter_4_11 ? hash_out_4_11 : 0;
    din_4_11.last <= out_new_pkt;
    din_4_11.bucket <= 4;


    din_4_11_r1 <= din_4_11;
    din_4_11_r2 <= din_4_11_r1;
    din_valid_4_12 <= out_new_pkt | hash_out_valid_filter_4_12;
    din_valid_4_12_r1 <= din_valid_4_12;
    din_valid_4_12_r2 <= din_valid_4_12_r1;

    din_4_12.data <= hash_out_valid_filter_4_12 ? hash_out_4_12 : 0;
    din_4_12.last <= out_new_pkt;
    din_4_12.bucket <= 4;


    din_4_12_r1 <= din_4_12;
    din_4_12_r2 <= din_4_12_r1;
    din_valid_4_13 <= out_new_pkt | hash_out_valid_filter_4_13;
    din_valid_4_13_r1 <= din_valid_4_13;
    din_valid_4_13_r2 <= din_valid_4_13_r1;

    din_4_13.data <= hash_out_valid_filter_4_13 ? hash_out_4_13 : 0;
    din_4_13.last <= out_new_pkt;
    din_4_13.bucket <= 4;


    din_4_13_r1 <= din_4_13;
    din_4_13_r2 <= din_4_13_r1;
    din_valid_4_14 <= out_new_pkt | hash_out_valid_filter_4_14;
    din_valid_4_14_r1 <= din_valid_4_14;
    din_valid_4_14_r2 <= din_valid_4_14_r1;

    din_4_14.data <= hash_out_valid_filter_4_14 ? hash_out_4_14 : 0;
    din_4_14.last <= out_new_pkt;
    din_4_14.bucket <= 4;


    din_4_14_r1 <= din_4_14;
    din_4_14_r2 <= din_4_14_r1;
    din_valid_4_15 <= out_new_pkt | hash_out_valid_filter_4_15;
    din_valid_4_15_r1 <= din_valid_4_15;
    din_valid_4_15_r2 <= din_valid_4_15_r1;

    din_4_15.data <= hash_out_valid_filter_4_15 ? hash_out_4_15 : 0;
    din_4_15.last <= out_new_pkt;
    din_4_15.bucket <= 4;


    din_4_15_r1 <= din_4_15;
    din_4_15_r2 <= din_4_15_r1;
    din_valid_4_16 <= out_new_pkt | hash_out_valid_filter_4_16;
    din_valid_4_16_r1 <= din_valid_4_16;
    din_valid_4_16_r2 <= din_valid_4_16_r1;

    din_4_16.data <= hash_out_valid_filter_4_16 ? hash_out_4_16 : 0;
    din_4_16.last <= out_new_pkt;
    din_4_16.bucket <= 4;


    din_4_16_r1 <= din_4_16;
    din_4_16_r2 <= din_4_16_r1;
    din_valid_4_17 <= out_new_pkt | hash_out_valid_filter_4_17;
    din_valid_4_17_r1 <= din_valid_4_17;
    din_valid_4_17_r2 <= din_valid_4_17_r1;

    din_4_17.data <= hash_out_valid_filter_4_17 ? hash_out_4_17 : 0;
    din_4_17.last <= out_new_pkt;
    din_4_17.bucket <= 4;


    din_4_17_r1 <= din_4_17;
    din_4_17_r2 <= din_4_17_r1;
    din_valid_4_18 <= out_new_pkt | hash_out_valid_filter_4_18;
    din_valid_4_18_r1 <= din_valid_4_18;
    din_valid_4_18_r2 <= din_valid_4_18_r1;

    din_4_18.data <= hash_out_valid_filter_4_18 ? hash_out_4_18 : 0;
    din_4_18.last <= out_new_pkt;
    din_4_18.bucket <= 4;


    din_4_18_r1 <= din_4_18;
    din_4_18_r2 <= din_4_18_r1;
    din_valid_4_19 <= out_new_pkt | hash_out_valid_filter_4_19;
    din_valid_4_19_r1 <= din_valid_4_19;
    din_valid_4_19_r2 <= din_valid_4_19_r1;

    din_4_19.data <= hash_out_valid_filter_4_19 ? hash_out_4_19 : 0;
    din_4_19.last <= out_new_pkt;
    din_4_19.bucket <= 4;


    din_4_19_r1 <= din_4_19;
    din_4_19_r2 <= din_4_19_r1;
    din_valid_4_20 <= out_new_pkt | hash_out_valid_filter_4_20;
    din_valid_4_20_r1 <= din_valid_4_20;
    din_valid_4_20_r2 <= din_valid_4_20_r1;

    din_4_20.data <= hash_out_valid_filter_4_20 ? hash_out_4_20 : 0;
    din_4_20.last <= out_new_pkt;
    din_4_20.bucket <= 4;


    din_4_20_r1 <= din_4_20;
    din_4_20_r2 <= din_4_20_r1;
    din_valid_4_21 <= out_new_pkt | hash_out_valid_filter_4_21;
    din_valid_4_21_r1 <= din_valid_4_21;
    din_valid_4_21_r2 <= din_valid_4_21_r1;

    din_4_21.data <= hash_out_valid_filter_4_21 ? hash_out_4_21 : 0;
    din_4_21.last <= out_new_pkt;
    din_4_21.bucket <= 4;


    din_4_21_r1 <= din_4_21;
    din_4_21_r2 <= din_4_21_r1;
    din_valid_4_22 <= out_new_pkt | hash_out_valid_filter_4_22;
    din_valid_4_22_r1 <= din_valid_4_22;
    din_valid_4_22_r2 <= din_valid_4_22_r1;

    din_4_22.data <= hash_out_valid_filter_4_22 ? hash_out_4_22 : 0;
    din_4_22.last <= out_new_pkt;
    din_4_22.bucket <= 4;


    din_4_22_r1 <= din_4_22;
    din_4_22_r2 <= din_4_22_r1;
    din_valid_4_23 <= out_new_pkt | hash_out_valid_filter_4_23;
    din_valid_4_23_r1 <= din_valid_4_23;
    din_valid_4_23_r2 <= din_valid_4_23_r1;

    din_4_23.data <= hash_out_valid_filter_4_23 ? hash_out_4_23 : 0;
    din_4_23.last <= out_new_pkt;
    din_4_23.bucket <= 4;


    din_4_23_r1 <= din_4_23;
    din_4_23_r2 <= din_4_23_r1;
    din_valid_4_24 <= out_new_pkt | hash_out_valid_filter_4_24;
    din_valid_4_24_r1 <= din_valid_4_24;
    din_valid_4_24_r2 <= din_valid_4_24_r1;

    din_4_24.data <= hash_out_valid_filter_4_24 ? hash_out_4_24 : 0;
    din_4_24.last <= out_new_pkt;
    din_4_24.bucket <= 4;


    din_4_24_r1 <= din_4_24;
    din_4_24_r2 <= din_4_24_r1;
    din_valid_4_25 <= out_new_pkt | hash_out_valid_filter_4_25;
    din_valid_4_25_r1 <= din_valid_4_25;
    din_valid_4_25_r2 <= din_valid_4_25_r1;

    din_4_25.data <= hash_out_valid_filter_4_25 ? hash_out_4_25 : 0;
    din_4_25.last <= out_new_pkt;
    din_4_25.bucket <= 4;


    din_4_25_r1 <= din_4_25;
    din_4_25_r2 <= din_4_25_r1;
    din_valid_4_26 <= out_new_pkt | hash_out_valid_filter_4_26;
    din_valid_4_26_r1 <= din_valid_4_26;
    din_valid_4_26_r2 <= din_valid_4_26_r1;

    din_4_26.data <= hash_out_valid_filter_4_26 ? hash_out_4_26 : 0;
    din_4_26.last <= out_new_pkt;
    din_4_26.bucket <= 4;


    din_4_26_r1 <= din_4_26;
    din_4_26_r2 <= din_4_26_r1;
    din_valid_4_27 <= out_new_pkt | hash_out_valid_filter_4_27;
    din_valid_4_27_r1 <= din_valid_4_27;
    din_valid_4_27_r2 <= din_valid_4_27_r1;

    din_4_27.data <= hash_out_valid_filter_4_27 ? hash_out_4_27 : 0;
    din_4_27.last <= out_new_pkt;
    din_4_27.bucket <= 4;


    din_4_27_r1 <= din_4_27;
    din_4_27_r2 <= din_4_27_r1;
    din_valid_4_28 <= out_new_pkt | hash_out_valid_filter_4_28;
    din_valid_4_28_r1 <= din_valid_4_28;
    din_valid_4_28_r2 <= din_valid_4_28_r1;

    din_4_28.data <= hash_out_valid_filter_4_28 ? hash_out_4_28 : 0;
    din_4_28.last <= out_new_pkt;
    din_4_28.bucket <= 4;


    din_4_28_r1 <= din_4_28;
    din_4_28_r2 <= din_4_28_r1;
    din_valid_4_29 <= out_new_pkt | hash_out_valid_filter_4_29;
    din_valid_4_29_r1 <= din_valid_4_29;
    din_valid_4_29_r2 <= din_valid_4_29_r1;

    din_4_29.data <= hash_out_valid_filter_4_29 ? hash_out_4_29 : 0;
    din_4_29.last <= out_new_pkt;
    din_4_29.bucket <= 4;


    din_4_29_r1 <= din_4_29;
    din_4_29_r2 <= din_4_29_r1;
    din_valid_4_30 <= out_new_pkt | hash_out_valid_filter_4_30;
    din_valid_4_30_r1 <= din_valid_4_30;
    din_valid_4_30_r2 <= din_valid_4_30_r1;

    din_4_30.data <= hash_out_valid_filter_4_30 ? hash_out_4_30 : 0;
    din_4_30.last <= out_new_pkt;
    din_4_30.bucket <= 4;


    din_4_30_r1 <= din_4_30;
    din_4_30_r2 <= din_4_30_r1;
    din_valid_4_31 <= out_new_pkt | hash_out_valid_filter_4_31;
    din_valid_4_31_r1 <= din_valid_4_31;
    din_valid_4_31_r2 <= din_valid_4_31_r1;

    din_4_31.data <= hash_out_valid_filter_4_31 ? hash_out_4_31 : 0;
    din_4_31.last <= out_new_pkt;
    din_4_31.bucket <= 4;


    din_4_31_r1 <= din_4_31;
    din_4_31_r2 <= din_4_31_r1;
    din_valid_5_0 <= out_new_pkt | hash_out_valid_filter_5_0;
    din_valid_5_0_r1 <= din_valid_5_0;
    din_valid_5_0_r2 <= din_valid_5_0_r1;

    din_5_0.data <= hash_out_valid_filter_5_0 ? hash_out_5_0 : 0;
    din_5_0.last <= out_new_pkt;
    din_5_0.bucket <= 5;


    din_5_0_r1 <= din_5_0;
    din_5_0_r2 <= din_5_0_r1;
    din_valid_5_1 <= out_new_pkt | hash_out_valid_filter_5_1;
    din_valid_5_1_r1 <= din_valid_5_1;
    din_valid_5_1_r2 <= din_valid_5_1_r1;

    din_5_1.data <= hash_out_valid_filter_5_1 ? hash_out_5_1 : 0;
    din_5_1.last <= out_new_pkt;
    din_5_1.bucket <= 5;


    din_5_1_r1 <= din_5_1;
    din_5_1_r2 <= din_5_1_r1;
    din_valid_5_2 <= out_new_pkt | hash_out_valid_filter_5_2;
    din_valid_5_2_r1 <= din_valid_5_2;
    din_valid_5_2_r2 <= din_valid_5_2_r1;

    din_5_2.data <= hash_out_valid_filter_5_2 ? hash_out_5_2 : 0;
    din_5_2.last <= out_new_pkt;
    din_5_2.bucket <= 5;


    din_5_2_r1 <= din_5_2;
    din_5_2_r2 <= din_5_2_r1;
    din_valid_5_3 <= out_new_pkt | hash_out_valid_filter_5_3;
    din_valid_5_3_r1 <= din_valid_5_3;
    din_valid_5_3_r2 <= din_valid_5_3_r1;

    din_5_3.data <= hash_out_valid_filter_5_3 ? hash_out_5_3 : 0;
    din_5_3.last <= out_new_pkt;
    din_5_3.bucket <= 5;


    din_5_3_r1 <= din_5_3;
    din_5_3_r2 <= din_5_3_r1;
    din_valid_5_4 <= out_new_pkt | hash_out_valid_filter_5_4;
    din_valid_5_4_r1 <= din_valid_5_4;
    din_valid_5_4_r2 <= din_valid_5_4_r1;

    din_5_4.data <= hash_out_valid_filter_5_4 ? hash_out_5_4 : 0;
    din_5_4.last <= out_new_pkt;
    din_5_4.bucket <= 5;


    din_5_4_r1 <= din_5_4;
    din_5_4_r2 <= din_5_4_r1;
    din_valid_5_5 <= out_new_pkt | hash_out_valid_filter_5_5;
    din_valid_5_5_r1 <= din_valid_5_5;
    din_valid_5_5_r2 <= din_valid_5_5_r1;

    din_5_5.data <= hash_out_valid_filter_5_5 ? hash_out_5_5 : 0;
    din_5_5.last <= out_new_pkt;
    din_5_5.bucket <= 5;


    din_5_5_r1 <= din_5_5;
    din_5_5_r2 <= din_5_5_r1;
    din_valid_5_6 <= out_new_pkt | hash_out_valid_filter_5_6;
    din_valid_5_6_r1 <= din_valid_5_6;
    din_valid_5_6_r2 <= din_valid_5_6_r1;

    din_5_6.data <= hash_out_valid_filter_5_6 ? hash_out_5_6 : 0;
    din_5_6.last <= out_new_pkt;
    din_5_6.bucket <= 5;


    din_5_6_r1 <= din_5_6;
    din_5_6_r2 <= din_5_6_r1;
    din_valid_5_7 <= out_new_pkt | hash_out_valid_filter_5_7;
    din_valid_5_7_r1 <= din_valid_5_7;
    din_valid_5_7_r2 <= din_valid_5_7_r1;

    din_5_7.data <= hash_out_valid_filter_5_7 ? hash_out_5_7 : 0;
    din_5_7.last <= out_new_pkt;
    din_5_7.bucket <= 5;


    din_5_7_r1 <= din_5_7;
    din_5_7_r2 <= din_5_7_r1;
    din_valid_5_8 <= out_new_pkt | hash_out_valid_filter_5_8;
    din_valid_5_8_r1 <= din_valid_5_8;
    din_valid_5_8_r2 <= din_valid_5_8_r1;

    din_5_8.data <= hash_out_valid_filter_5_8 ? hash_out_5_8 : 0;
    din_5_8.last <= out_new_pkt;
    din_5_8.bucket <= 5;


    din_5_8_r1 <= din_5_8;
    din_5_8_r2 <= din_5_8_r1;
    din_valid_5_9 <= out_new_pkt | hash_out_valid_filter_5_9;
    din_valid_5_9_r1 <= din_valid_5_9;
    din_valid_5_9_r2 <= din_valid_5_9_r1;

    din_5_9.data <= hash_out_valid_filter_5_9 ? hash_out_5_9 : 0;
    din_5_9.last <= out_new_pkt;
    din_5_9.bucket <= 5;


    din_5_9_r1 <= din_5_9;
    din_5_9_r2 <= din_5_9_r1;
    din_valid_5_10 <= out_new_pkt | hash_out_valid_filter_5_10;
    din_valid_5_10_r1 <= din_valid_5_10;
    din_valid_5_10_r2 <= din_valid_5_10_r1;

    din_5_10.data <= hash_out_valid_filter_5_10 ? hash_out_5_10 : 0;
    din_5_10.last <= out_new_pkt;
    din_5_10.bucket <= 5;


    din_5_10_r1 <= din_5_10;
    din_5_10_r2 <= din_5_10_r1;
    din_valid_5_11 <= out_new_pkt | hash_out_valid_filter_5_11;
    din_valid_5_11_r1 <= din_valid_5_11;
    din_valid_5_11_r2 <= din_valid_5_11_r1;

    din_5_11.data <= hash_out_valid_filter_5_11 ? hash_out_5_11 : 0;
    din_5_11.last <= out_new_pkt;
    din_5_11.bucket <= 5;


    din_5_11_r1 <= din_5_11;
    din_5_11_r2 <= din_5_11_r1;
    din_valid_5_12 <= out_new_pkt | hash_out_valid_filter_5_12;
    din_valid_5_12_r1 <= din_valid_5_12;
    din_valid_5_12_r2 <= din_valid_5_12_r1;

    din_5_12.data <= hash_out_valid_filter_5_12 ? hash_out_5_12 : 0;
    din_5_12.last <= out_new_pkt;
    din_5_12.bucket <= 5;


    din_5_12_r1 <= din_5_12;
    din_5_12_r2 <= din_5_12_r1;
    din_valid_5_13 <= out_new_pkt | hash_out_valid_filter_5_13;
    din_valid_5_13_r1 <= din_valid_5_13;
    din_valid_5_13_r2 <= din_valid_5_13_r1;

    din_5_13.data <= hash_out_valid_filter_5_13 ? hash_out_5_13 : 0;
    din_5_13.last <= out_new_pkt;
    din_5_13.bucket <= 5;


    din_5_13_r1 <= din_5_13;
    din_5_13_r2 <= din_5_13_r1;
    din_valid_5_14 <= out_new_pkt | hash_out_valid_filter_5_14;
    din_valid_5_14_r1 <= din_valid_5_14;
    din_valid_5_14_r2 <= din_valid_5_14_r1;

    din_5_14.data <= hash_out_valid_filter_5_14 ? hash_out_5_14 : 0;
    din_5_14.last <= out_new_pkt;
    din_5_14.bucket <= 5;


    din_5_14_r1 <= din_5_14;
    din_5_14_r2 <= din_5_14_r1;
    din_valid_5_15 <= out_new_pkt | hash_out_valid_filter_5_15;
    din_valid_5_15_r1 <= din_valid_5_15;
    din_valid_5_15_r2 <= din_valid_5_15_r1;

    din_5_15.data <= hash_out_valid_filter_5_15 ? hash_out_5_15 : 0;
    din_5_15.last <= out_new_pkt;
    din_5_15.bucket <= 5;


    din_5_15_r1 <= din_5_15;
    din_5_15_r2 <= din_5_15_r1;
    din_valid_5_16 <= out_new_pkt | hash_out_valid_filter_5_16;
    din_valid_5_16_r1 <= din_valid_5_16;
    din_valid_5_16_r2 <= din_valid_5_16_r1;

    din_5_16.data <= hash_out_valid_filter_5_16 ? hash_out_5_16 : 0;
    din_5_16.last <= out_new_pkt;
    din_5_16.bucket <= 5;


    din_5_16_r1 <= din_5_16;
    din_5_16_r2 <= din_5_16_r1;
    din_valid_5_17 <= out_new_pkt | hash_out_valid_filter_5_17;
    din_valid_5_17_r1 <= din_valid_5_17;
    din_valid_5_17_r2 <= din_valid_5_17_r1;

    din_5_17.data <= hash_out_valid_filter_5_17 ? hash_out_5_17 : 0;
    din_5_17.last <= out_new_pkt;
    din_5_17.bucket <= 5;


    din_5_17_r1 <= din_5_17;
    din_5_17_r2 <= din_5_17_r1;
    din_valid_5_18 <= out_new_pkt | hash_out_valid_filter_5_18;
    din_valid_5_18_r1 <= din_valid_5_18;
    din_valid_5_18_r2 <= din_valid_5_18_r1;

    din_5_18.data <= hash_out_valid_filter_5_18 ? hash_out_5_18 : 0;
    din_5_18.last <= out_new_pkt;
    din_5_18.bucket <= 5;


    din_5_18_r1 <= din_5_18;
    din_5_18_r2 <= din_5_18_r1;
    din_valid_5_19 <= out_new_pkt | hash_out_valid_filter_5_19;
    din_valid_5_19_r1 <= din_valid_5_19;
    din_valid_5_19_r2 <= din_valid_5_19_r1;

    din_5_19.data <= hash_out_valid_filter_5_19 ? hash_out_5_19 : 0;
    din_5_19.last <= out_new_pkt;
    din_5_19.bucket <= 5;


    din_5_19_r1 <= din_5_19;
    din_5_19_r2 <= din_5_19_r1;
    din_valid_5_20 <= out_new_pkt | hash_out_valid_filter_5_20;
    din_valid_5_20_r1 <= din_valid_5_20;
    din_valid_5_20_r2 <= din_valid_5_20_r1;

    din_5_20.data <= hash_out_valid_filter_5_20 ? hash_out_5_20 : 0;
    din_5_20.last <= out_new_pkt;
    din_5_20.bucket <= 5;


    din_5_20_r1 <= din_5_20;
    din_5_20_r2 <= din_5_20_r1;
    din_valid_5_21 <= out_new_pkt | hash_out_valid_filter_5_21;
    din_valid_5_21_r1 <= din_valid_5_21;
    din_valid_5_21_r2 <= din_valid_5_21_r1;

    din_5_21.data <= hash_out_valid_filter_5_21 ? hash_out_5_21 : 0;
    din_5_21.last <= out_new_pkt;
    din_5_21.bucket <= 5;


    din_5_21_r1 <= din_5_21;
    din_5_21_r2 <= din_5_21_r1;
    din_valid_5_22 <= out_new_pkt | hash_out_valid_filter_5_22;
    din_valid_5_22_r1 <= din_valid_5_22;
    din_valid_5_22_r2 <= din_valid_5_22_r1;

    din_5_22.data <= hash_out_valid_filter_5_22 ? hash_out_5_22 : 0;
    din_5_22.last <= out_new_pkt;
    din_5_22.bucket <= 5;


    din_5_22_r1 <= din_5_22;
    din_5_22_r2 <= din_5_22_r1;
    din_valid_5_23 <= out_new_pkt | hash_out_valid_filter_5_23;
    din_valid_5_23_r1 <= din_valid_5_23;
    din_valid_5_23_r2 <= din_valid_5_23_r1;

    din_5_23.data <= hash_out_valid_filter_5_23 ? hash_out_5_23 : 0;
    din_5_23.last <= out_new_pkt;
    din_5_23.bucket <= 5;


    din_5_23_r1 <= din_5_23;
    din_5_23_r2 <= din_5_23_r1;
    din_valid_5_24 <= out_new_pkt | hash_out_valid_filter_5_24;
    din_valid_5_24_r1 <= din_valid_5_24;
    din_valid_5_24_r2 <= din_valid_5_24_r1;

    din_5_24.data <= hash_out_valid_filter_5_24 ? hash_out_5_24 : 0;
    din_5_24.last <= out_new_pkt;
    din_5_24.bucket <= 5;


    din_5_24_r1 <= din_5_24;
    din_5_24_r2 <= din_5_24_r1;
    din_valid_5_25 <= out_new_pkt | hash_out_valid_filter_5_25;
    din_valid_5_25_r1 <= din_valid_5_25;
    din_valid_5_25_r2 <= din_valid_5_25_r1;

    din_5_25.data <= hash_out_valid_filter_5_25 ? hash_out_5_25 : 0;
    din_5_25.last <= out_new_pkt;
    din_5_25.bucket <= 5;


    din_5_25_r1 <= din_5_25;
    din_5_25_r2 <= din_5_25_r1;
    din_valid_5_26 <= out_new_pkt | hash_out_valid_filter_5_26;
    din_valid_5_26_r1 <= din_valid_5_26;
    din_valid_5_26_r2 <= din_valid_5_26_r1;

    din_5_26.data <= hash_out_valid_filter_5_26 ? hash_out_5_26 : 0;
    din_5_26.last <= out_new_pkt;
    din_5_26.bucket <= 5;


    din_5_26_r1 <= din_5_26;
    din_5_26_r2 <= din_5_26_r1;
    din_valid_5_27 <= out_new_pkt | hash_out_valid_filter_5_27;
    din_valid_5_27_r1 <= din_valid_5_27;
    din_valid_5_27_r2 <= din_valid_5_27_r1;

    din_5_27.data <= hash_out_valid_filter_5_27 ? hash_out_5_27 : 0;
    din_5_27.last <= out_new_pkt;
    din_5_27.bucket <= 5;


    din_5_27_r1 <= din_5_27;
    din_5_27_r2 <= din_5_27_r1;
    din_valid_5_28 <= out_new_pkt | hash_out_valid_filter_5_28;
    din_valid_5_28_r1 <= din_valid_5_28;
    din_valid_5_28_r2 <= din_valid_5_28_r1;

    din_5_28.data <= hash_out_valid_filter_5_28 ? hash_out_5_28 : 0;
    din_5_28.last <= out_new_pkt;
    din_5_28.bucket <= 5;


    din_5_28_r1 <= din_5_28;
    din_5_28_r2 <= din_5_28_r1;
    din_valid_5_29 <= out_new_pkt | hash_out_valid_filter_5_29;
    din_valid_5_29_r1 <= din_valid_5_29;
    din_valid_5_29_r2 <= din_valid_5_29_r1;

    din_5_29.data <= hash_out_valid_filter_5_29 ? hash_out_5_29 : 0;
    din_5_29.last <= out_new_pkt;
    din_5_29.bucket <= 5;


    din_5_29_r1 <= din_5_29;
    din_5_29_r2 <= din_5_29_r1;
    din_valid_5_30 <= out_new_pkt | hash_out_valid_filter_5_30;
    din_valid_5_30_r1 <= din_valid_5_30;
    din_valid_5_30_r2 <= din_valid_5_30_r1;

    din_5_30.data <= hash_out_valid_filter_5_30 ? hash_out_5_30 : 0;
    din_5_30.last <= out_new_pkt;
    din_5_30.bucket <= 5;


    din_5_30_r1 <= din_5_30;
    din_5_30_r2 <= din_5_30_r1;
    din_valid_5_31 <= out_new_pkt | hash_out_valid_filter_5_31;
    din_valid_5_31_r1 <= din_valid_5_31;
    din_valid_5_31_r2 <= din_valid_5_31_r1;

    din_5_31.data <= hash_out_valid_filter_5_31 ? hash_out_5_31 : 0;
    din_5_31.last <= out_new_pkt;
    din_5_31.bucket <= 5;


    din_5_31_r1 <= din_5_31;
    din_5_31_r2 <= din_5_31_r1;
    din_valid_6_0 <= out_new_pkt | hash_out_valid_filter_6_0;
    din_valid_6_0_r1 <= din_valid_6_0;
    din_valid_6_0_r2 <= din_valid_6_0_r1;

    din_6_0.data <= hash_out_valid_filter_6_0 ? hash_out_6_0 : 0;
    din_6_0.last <= out_new_pkt;
    din_6_0.bucket <= 6;


    din_6_0_r1 <= din_6_0;
    din_6_0_r2 <= din_6_0_r1;
    din_valid_6_1 <= out_new_pkt | hash_out_valid_filter_6_1;
    din_valid_6_1_r1 <= din_valid_6_1;
    din_valid_6_1_r2 <= din_valid_6_1_r1;

    din_6_1.data <= hash_out_valid_filter_6_1 ? hash_out_6_1 : 0;
    din_6_1.last <= out_new_pkt;
    din_6_1.bucket <= 6;


    din_6_1_r1 <= din_6_1;
    din_6_1_r2 <= din_6_1_r1;
    din_valid_6_2 <= out_new_pkt | hash_out_valid_filter_6_2;
    din_valid_6_2_r1 <= din_valid_6_2;
    din_valid_6_2_r2 <= din_valid_6_2_r1;

    din_6_2.data <= hash_out_valid_filter_6_2 ? hash_out_6_2 : 0;
    din_6_2.last <= out_new_pkt;
    din_6_2.bucket <= 6;


    din_6_2_r1 <= din_6_2;
    din_6_2_r2 <= din_6_2_r1;
    din_valid_6_3 <= out_new_pkt | hash_out_valid_filter_6_3;
    din_valid_6_3_r1 <= din_valid_6_3;
    din_valid_6_3_r2 <= din_valid_6_3_r1;

    din_6_3.data <= hash_out_valid_filter_6_3 ? hash_out_6_3 : 0;
    din_6_3.last <= out_new_pkt;
    din_6_3.bucket <= 6;


    din_6_3_r1 <= din_6_3;
    din_6_3_r2 <= din_6_3_r1;
    din_valid_6_4 <= out_new_pkt | hash_out_valid_filter_6_4;
    din_valid_6_4_r1 <= din_valid_6_4;
    din_valid_6_4_r2 <= din_valid_6_4_r1;

    din_6_4.data <= hash_out_valid_filter_6_4 ? hash_out_6_4 : 0;
    din_6_4.last <= out_new_pkt;
    din_6_4.bucket <= 6;


    din_6_4_r1 <= din_6_4;
    din_6_4_r2 <= din_6_4_r1;
    din_valid_6_5 <= out_new_pkt | hash_out_valid_filter_6_5;
    din_valid_6_5_r1 <= din_valid_6_5;
    din_valid_6_5_r2 <= din_valid_6_5_r1;

    din_6_5.data <= hash_out_valid_filter_6_5 ? hash_out_6_5 : 0;
    din_6_5.last <= out_new_pkt;
    din_6_5.bucket <= 6;


    din_6_5_r1 <= din_6_5;
    din_6_5_r2 <= din_6_5_r1;
    din_valid_6_6 <= out_new_pkt | hash_out_valid_filter_6_6;
    din_valid_6_6_r1 <= din_valid_6_6;
    din_valid_6_6_r2 <= din_valid_6_6_r1;

    din_6_6.data <= hash_out_valid_filter_6_6 ? hash_out_6_6 : 0;
    din_6_6.last <= out_new_pkt;
    din_6_6.bucket <= 6;


    din_6_6_r1 <= din_6_6;
    din_6_6_r2 <= din_6_6_r1;
    din_valid_6_7 <= out_new_pkt | hash_out_valid_filter_6_7;
    din_valid_6_7_r1 <= din_valid_6_7;
    din_valid_6_7_r2 <= din_valid_6_7_r1;

    din_6_7.data <= hash_out_valid_filter_6_7 ? hash_out_6_7 : 0;
    din_6_7.last <= out_new_pkt;
    din_6_7.bucket <= 6;


    din_6_7_r1 <= din_6_7;
    din_6_7_r2 <= din_6_7_r1;
    din_valid_6_8 <= out_new_pkt | hash_out_valid_filter_6_8;
    din_valid_6_8_r1 <= din_valid_6_8;
    din_valid_6_8_r2 <= din_valid_6_8_r1;

    din_6_8.data <= hash_out_valid_filter_6_8 ? hash_out_6_8 : 0;
    din_6_8.last <= out_new_pkt;
    din_6_8.bucket <= 6;


    din_6_8_r1 <= din_6_8;
    din_6_8_r2 <= din_6_8_r1;
    din_valid_6_9 <= out_new_pkt | hash_out_valid_filter_6_9;
    din_valid_6_9_r1 <= din_valid_6_9;
    din_valid_6_9_r2 <= din_valid_6_9_r1;

    din_6_9.data <= hash_out_valid_filter_6_9 ? hash_out_6_9 : 0;
    din_6_9.last <= out_new_pkt;
    din_6_9.bucket <= 6;


    din_6_9_r1 <= din_6_9;
    din_6_9_r2 <= din_6_9_r1;
    din_valid_6_10 <= out_new_pkt | hash_out_valid_filter_6_10;
    din_valid_6_10_r1 <= din_valid_6_10;
    din_valid_6_10_r2 <= din_valid_6_10_r1;

    din_6_10.data <= hash_out_valid_filter_6_10 ? hash_out_6_10 : 0;
    din_6_10.last <= out_new_pkt;
    din_6_10.bucket <= 6;


    din_6_10_r1 <= din_6_10;
    din_6_10_r2 <= din_6_10_r1;
    din_valid_6_11 <= out_new_pkt | hash_out_valid_filter_6_11;
    din_valid_6_11_r1 <= din_valid_6_11;
    din_valid_6_11_r2 <= din_valid_6_11_r1;

    din_6_11.data <= hash_out_valid_filter_6_11 ? hash_out_6_11 : 0;
    din_6_11.last <= out_new_pkt;
    din_6_11.bucket <= 6;


    din_6_11_r1 <= din_6_11;
    din_6_11_r2 <= din_6_11_r1;
    din_valid_6_12 <= out_new_pkt | hash_out_valid_filter_6_12;
    din_valid_6_12_r1 <= din_valid_6_12;
    din_valid_6_12_r2 <= din_valid_6_12_r1;

    din_6_12.data <= hash_out_valid_filter_6_12 ? hash_out_6_12 : 0;
    din_6_12.last <= out_new_pkt;
    din_6_12.bucket <= 6;


    din_6_12_r1 <= din_6_12;
    din_6_12_r2 <= din_6_12_r1;
    din_valid_6_13 <= out_new_pkt | hash_out_valid_filter_6_13;
    din_valid_6_13_r1 <= din_valid_6_13;
    din_valid_6_13_r2 <= din_valid_6_13_r1;

    din_6_13.data <= hash_out_valid_filter_6_13 ? hash_out_6_13 : 0;
    din_6_13.last <= out_new_pkt;
    din_6_13.bucket <= 6;


    din_6_13_r1 <= din_6_13;
    din_6_13_r2 <= din_6_13_r1;
    din_valid_6_14 <= out_new_pkt | hash_out_valid_filter_6_14;
    din_valid_6_14_r1 <= din_valid_6_14;
    din_valid_6_14_r2 <= din_valid_6_14_r1;

    din_6_14.data <= hash_out_valid_filter_6_14 ? hash_out_6_14 : 0;
    din_6_14.last <= out_new_pkt;
    din_6_14.bucket <= 6;


    din_6_14_r1 <= din_6_14;
    din_6_14_r2 <= din_6_14_r1;
    din_valid_6_15 <= out_new_pkt | hash_out_valid_filter_6_15;
    din_valid_6_15_r1 <= din_valid_6_15;
    din_valid_6_15_r2 <= din_valid_6_15_r1;

    din_6_15.data <= hash_out_valid_filter_6_15 ? hash_out_6_15 : 0;
    din_6_15.last <= out_new_pkt;
    din_6_15.bucket <= 6;


    din_6_15_r1 <= din_6_15;
    din_6_15_r2 <= din_6_15_r1;
    din_valid_6_16 <= out_new_pkt | hash_out_valid_filter_6_16;
    din_valid_6_16_r1 <= din_valid_6_16;
    din_valid_6_16_r2 <= din_valid_6_16_r1;

    din_6_16.data <= hash_out_valid_filter_6_16 ? hash_out_6_16 : 0;
    din_6_16.last <= out_new_pkt;
    din_6_16.bucket <= 6;


    din_6_16_r1 <= din_6_16;
    din_6_16_r2 <= din_6_16_r1;
    din_valid_6_17 <= out_new_pkt | hash_out_valid_filter_6_17;
    din_valid_6_17_r1 <= din_valid_6_17;
    din_valid_6_17_r2 <= din_valid_6_17_r1;

    din_6_17.data <= hash_out_valid_filter_6_17 ? hash_out_6_17 : 0;
    din_6_17.last <= out_new_pkt;
    din_6_17.bucket <= 6;


    din_6_17_r1 <= din_6_17;
    din_6_17_r2 <= din_6_17_r1;
    din_valid_6_18 <= out_new_pkt | hash_out_valid_filter_6_18;
    din_valid_6_18_r1 <= din_valid_6_18;
    din_valid_6_18_r2 <= din_valid_6_18_r1;

    din_6_18.data <= hash_out_valid_filter_6_18 ? hash_out_6_18 : 0;
    din_6_18.last <= out_new_pkt;
    din_6_18.bucket <= 6;


    din_6_18_r1 <= din_6_18;
    din_6_18_r2 <= din_6_18_r1;
    din_valid_6_19 <= out_new_pkt | hash_out_valid_filter_6_19;
    din_valid_6_19_r1 <= din_valid_6_19;
    din_valid_6_19_r2 <= din_valid_6_19_r1;

    din_6_19.data <= hash_out_valid_filter_6_19 ? hash_out_6_19 : 0;
    din_6_19.last <= out_new_pkt;
    din_6_19.bucket <= 6;


    din_6_19_r1 <= din_6_19;
    din_6_19_r2 <= din_6_19_r1;
    din_valid_6_20 <= out_new_pkt | hash_out_valid_filter_6_20;
    din_valid_6_20_r1 <= din_valid_6_20;
    din_valid_6_20_r2 <= din_valid_6_20_r1;

    din_6_20.data <= hash_out_valid_filter_6_20 ? hash_out_6_20 : 0;
    din_6_20.last <= out_new_pkt;
    din_6_20.bucket <= 6;


    din_6_20_r1 <= din_6_20;
    din_6_20_r2 <= din_6_20_r1;
    din_valid_6_21 <= out_new_pkt | hash_out_valid_filter_6_21;
    din_valid_6_21_r1 <= din_valid_6_21;
    din_valid_6_21_r2 <= din_valid_6_21_r1;

    din_6_21.data <= hash_out_valid_filter_6_21 ? hash_out_6_21 : 0;
    din_6_21.last <= out_new_pkt;
    din_6_21.bucket <= 6;


    din_6_21_r1 <= din_6_21;
    din_6_21_r2 <= din_6_21_r1;
    din_valid_6_22 <= out_new_pkt | hash_out_valid_filter_6_22;
    din_valid_6_22_r1 <= din_valid_6_22;
    din_valid_6_22_r2 <= din_valid_6_22_r1;

    din_6_22.data <= hash_out_valid_filter_6_22 ? hash_out_6_22 : 0;
    din_6_22.last <= out_new_pkt;
    din_6_22.bucket <= 6;


    din_6_22_r1 <= din_6_22;
    din_6_22_r2 <= din_6_22_r1;
    din_valid_6_23 <= out_new_pkt | hash_out_valid_filter_6_23;
    din_valid_6_23_r1 <= din_valid_6_23;
    din_valid_6_23_r2 <= din_valid_6_23_r1;

    din_6_23.data <= hash_out_valid_filter_6_23 ? hash_out_6_23 : 0;
    din_6_23.last <= out_new_pkt;
    din_6_23.bucket <= 6;


    din_6_23_r1 <= din_6_23;
    din_6_23_r2 <= din_6_23_r1;
    din_valid_6_24 <= out_new_pkt | hash_out_valid_filter_6_24;
    din_valid_6_24_r1 <= din_valid_6_24;
    din_valid_6_24_r2 <= din_valid_6_24_r1;

    din_6_24.data <= hash_out_valid_filter_6_24 ? hash_out_6_24 : 0;
    din_6_24.last <= out_new_pkt;
    din_6_24.bucket <= 6;


    din_6_24_r1 <= din_6_24;
    din_6_24_r2 <= din_6_24_r1;
    din_valid_6_25 <= out_new_pkt | hash_out_valid_filter_6_25;
    din_valid_6_25_r1 <= din_valid_6_25;
    din_valid_6_25_r2 <= din_valid_6_25_r1;

    din_6_25.data <= hash_out_valid_filter_6_25 ? hash_out_6_25 : 0;
    din_6_25.last <= out_new_pkt;
    din_6_25.bucket <= 6;


    din_6_25_r1 <= din_6_25;
    din_6_25_r2 <= din_6_25_r1;
    din_valid_6_26 <= out_new_pkt | hash_out_valid_filter_6_26;
    din_valid_6_26_r1 <= din_valid_6_26;
    din_valid_6_26_r2 <= din_valid_6_26_r1;

    din_6_26.data <= hash_out_valid_filter_6_26 ? hash_out_6_26 : 0;
    din_6_26.last <= out_new_pkt;
    din_6_26.bucket <= 6;


    din_6_26_r1 <= din_6_26;
    din_6_26_r2 <= din_6_26_r1;
    din_valid_6_27 <= out_new_pkt | hash_out_valid_filter_6_27;
    din_valid_6_27_r1 <= din_valid_6_27;
    din_valid_6_27_r2 <= din_valid_6_27_r1;

    din_6_27.data <= hash_out_valid_filter_6_27 ? hash_out_6_27 : 0;
    din_6_27.last <= out_new_pkt;
    din_6_27.bucket <= 6;


    din_6_27_r1 <= din_6_27;
    din_6_27_r2 <= din_6_27_r1;
    din_valid_6_28 <= out_new_pkt | hash_out_valid_filter_6_28;
    din_valid_6_28_r1 <= din_valid_6_28;
    din_valid_6_28_r2 <= din_valid_6_28_r1;

    din_6_28.data <= hash_out_valid_filter_6_28 ? hash_out_6_28 : 0;
    din_6_28.last <= out_new_pkt;
    din_6_28.bucket <= 6;


    din_6_28_r1 <= din_6_28;
    din_6_28_r2 <= din_6_28_r1;
    din_valid_6_29 <= out_new_pkt | hash_out_valid_filter_6_29;
    din_valid_6_29_r1 <= din_valid_6_29;
    din_valid_6_29_r2 <= din_valid_6_29_r1;

    din_6_29.data <= hash_out_valid_filter_6_29 ? hash_out_6_29 : 0;
    din_6_29.last <= out_new_pkt;
    din_6_29.bucket <= 6;


    din_6_29_r1 <= din_6_29;
    din_6_29_r2 <= din_6_29_r1;
    din_valid_6_30 <= out_new_pkt | hash_out_valid_filter_6_30;
    din_valid_6_30_r1 <= din_valid_6_30;
    din_valid_6_30_r2 <= din_valid_6_30_r1;

    din_6_30.data <= hash_out_valid_filter_6_30 ? hash_out_6_30 : 0;
    din_6_30.last <= out_new_pkt;
    din_6_30.bucket <= 6;


    din_6_30_r1 <= din_6_30;
    din_6_30_r2 <= din_6_30_r1;
    din_valid_6_31 <= out_new_pkt | hash_out_valid_filter_6_31;
    din_valid_6_31_r1 <= din_valid_6_31;
    din_valid_6_31_r2 <= din_valid_6_31_r1;

    din_6_31.data <= hash_out_valid_filter_6_31 ? hash_out_6_31 : 0;
    din_6_31.last <= out_new_pkt;
    din_6_31.bucket <= 6;


    din_6_31_r1 <= din_6_31;
    din_6_31_r2 <= din_6_31_r1;
    din_valid_7_0 <= out_new_pkt | hash_out_valid_filter_7_0;
    din_valid_7_0_r1 <= din_valid_7_0;
    din_valid_7_0_r2 <= din_valid_7_0_r1;

    din_7_0.data <= hash_out_valid_filter_7_0 ? hash_out_7_0 : 0;
    din_7_0.last <= out_new_pkt;
    din_7_0.bucket <= 7;


    din_7_0_r1 <= din_7_0;
    din_7_0_r2 <= din_7_0_r1;
    din_valid_7_1 <= out_new_pkt | hash_out_valid_filter_7_1;
    din_valid_7_1_r1 <= din_valid_7_1;
    din_valid_7_1_r2 <= din_valid_7_1_r1;

    din_7_1.data <= hash_out_valid_filter_7_1 ? hash_out_7_1 : 0;
    din_7_1.last <= out_new_pkt;
    din_7_1.bucket <= 7;


    din_7_1_r1 <= din_7_1;
    din_7_1_r2 <= din_7_1_r1;
    din_valid_7_2 <= out_new_pkt | hash_out_valid_filter_7_2;
    din_valid_7_2_r1 <= din_valid_7_2;
    din_valid_7_2_r2 <= din_valid_7_2_r1;

    din_7_2.data <= hash_out_valid_filter_7_2 ? hash_out_7_2 : 0;
    din_7_2.last <= out_new_pkt;
    din_7_2.bucket <= 7;


    din_7_2_r1 <= din_7_2;
    din_7_2_r2 <= din_7_2_r1;
    din_valid_7_3 <= out_new_pkt | hash_out_valid_filter_7_3;
    din_valid_7_3_r1 <= din_valid_7_3;
    din_valid_7_3_r2 <= din_valid_7_3_r1;

    din_7_3.data <= hash_out_valid_filter_7_3 ? hash_out_7_3 : 0;
    din_7_3.last <= out_new_pkt;
    din_7_3.bucket <= 7;


    din_7_3_r1 <= din_7_3;
    din_7_3_r2 <= din_7_3_r1;
    din_valid_7_4 <= out_new_pkt | hash_out_valid_filter_7_4;
    din_valid_7_4_r1 <= din_valid_7_4;
    din_valid_7_4_r2 <= din_valid_7_4_r1;

    din_7_4.data <= hash_out_valid_filter_7_4 ? hash_out_7_4 : 0;
    din_7_4.last <= out_new_pkt;
    din_7_4.bucket <= 7;


    din_7_4_r1 <= din_7_4;
    din_7_4_r2 <= din_7_4_r1;
    din_valid_7_5 <= out_new_pkt | hash_out_valid_filter_7_5;
    din_valid_7_5_r1 <= din_valid_7_5;
    din_valid_7_5_r2 <= din_valid_7_5_r1;

    din_7_5.data <= hash_out_valid_filter_7_5 ? hash_out_7_5 : 0;
    din_7_5.last <= out_new_pkt;
    din_7_5.bucket <= 7;


    din_7_5_r1 <= din_7_5;
    din_7_5_r2 <= din_7_5_r1;
    din_valid_7_6 <= out_new_pkt | hash_out_valid_filter_7_6;
    din_valid_7_6_r1 <= din_valid_7_6;
    din_valid_7_6_r2 <= din_valid_7_6_r1;

    din_7_6.data <= hash_out_valid_filter_7_6 ? hash_out_7_6 : 0;
    din_7_6.last <= out_new_pkt;
    din_7_6.bucket <= 7;


    din_7_6_r1 <= din_7_6;
    din_7_6_r2 <= din_7_6_r1;
    din_valid_7_7 <= out_new_pkt | hash_out_valid_filter_7_7;
    din_valid_7_7_r1 <= din_valid_7_7;
    din_valid_7_7_r2 <= din_valid_7_7_r1;

    din_7_7.data <= hash_out_valid_filter_7_7 ? hash_out_7_7 : 0;
    din_7_7.last <= out_new_pkt;
    din_7_7.bucket <= 7;


    din_7_7_r1 <= din_7_7;
    din_7_7_r2 <= din_7_7_r1;
    din_valid_7_8 <= out_new_pkt | hash_out_valid_filter_7_8;
    din_valid_7_8_r1 <= din_valid_7_8;
    din_valid_7_8_r2 <= din_valid_7_8_r1;

    din_7_8.data <= hash_out_valid_filter_7_8 ? hash_out_7_8 : 0;
    din_7_8.last <= out_new_pkt;
    din_7_8.bucket <= 7;


    din_7_8_r1 <= din_7_8;
    din_7_8_r2 <= din_7_8_r1;
    din_valid_7_9 <= out_new_pkt | hash_out_valid_filter_7_9;
    din_valid_7_9_r1 <= din_valid_7_9;
    din_valid_7_9_r2 <= din_valid_7_9_r1;

    din_7_9.data <= hash_out_valid_filter_7_9 ? hash_out_7_9 : 0;
    din_7_9.last <= out_new_pkt;
    din_7_9.bucket <= 7;


    din_7_9_r1 <= din_7_9;
    din_7_9_r2 <= din_7_9_r1;
    din_valid_7_10 <= out_new_pkt | hash_out_valid_filter_7_10;
    din_valid_7_10_r1 <= din_valid_7_10;
    din_valid_7_10_r2 <= din_valid_7_10_r1;

    din_7_10.data <= hash_out_valid_filter_7_10 ? hash_out_7_10 : 0;
    din_7_10.last <= out_new_pkt;
    din_7_10.bucket <= 7;


    din_7_10_r1 <= din_7_10;
    din_7_10_r2 <= din_7_10_r1;
    din_valid_7_11 <= out_new_pkt | hash_out_valid_filter_7_11;
    din_valid_7_11_r1 <= din_valid_7_11;
    din_valid_7_11_r2 <= din_valid_7_11_r1;

    din_7_11.data <= hash_out_valid_filter_7_11 ? hash_out_7_11 : 0;
    din_7_11.last <= out_new_pkt;
    din_7_11.bucket <= 7;


    din_7_11_r1 <= din_7_11;
    din_7_11_r2 <= din_7_11_r1;
    din_valid_7_12 <= out_new_pkt | hash_out_valid_filter_7_12;
    din_valid_7_12_r1 <= din_valid_7_12;
    din_valid_7_12_r2 <= din_valid_7_12_r1;

    din_7_12.data <= hash_out_valid_filter_7_12 ? hash_out_7_12 : 0;
    din_7_12.last <= out_new_pkt;
    din_7_12.bucket <= 7;


    din_7_12_r1 <= din_7_12;
    din_7_12_r2 <= din_7_12_r1;
    din_valid_7_13 <= out_new_pkt | hash_out_valid_filter_7_13;
    din_valid_7_13_r1 <= din_valid_7_13;
    din_valid_7_13_r2 <= din_valid_7_13_r1;

    din_7_13.data <= hash_out_valid_filter_7_13 ? hash_out_7_13 : 0;
    din_7_13.last <= out_new_pkt;
    din_7_13.bucket <= 7;


    din_7_13_r1 <= din_7_13;
    din_7_13_r2 <= din_7_13_r1;
    din_valid_7_14 <= out_new_pkt | hash_out_valid_filter_7_14;
    din_valid_7_14_r1 <= din_valid_7_14;
    din_valid_7_14_r2 <= din_valid_7_14_r1;

    din_7_14.data <= hash_out_valid_filter_7_14 ? hash_out_7_14 : 0;
    din_7_14.last <= out_new_pkt;
    din_7_14.bucket <= 7;


    din_7_14_r1 <= din_7_14;
    din_7_14_r2 <= din_7_14_r1;
    din_valid_7_15 <= out_new_pkt | hash_out_valid_filter_7_15;
    din_valid_7_15_r1 <= din_valid_7_15;
    din_valid_7_15_r2 <= din_valid_7_15_r1;

    din_7_15.data <= hash_out_valid_filter_7_15 ? hash_out_7_15 : 0;
    din_7_15.last <= out_new_pkt;
    din_7_15.bucket <= 7;


    din_7_15_r1 <= din_7_15;
    din_7_15_r2 <= din_7_15_r1;
    din_valid_7_16 <= out_new_pkt | hash_out_valid_filter_7_16;
    din_valid_7_16_r1 <= din_valid_7_16;
    din_valid_7_16_r2 <= din_valid_7_16_r1;

    din_7_16.data <= hash_out_valid_filter_7_16 ? hash_out_7_16 : 0;
    din_7_16.last <= out_new_pkt;
    din_7_16.bucket <= 7;


    din_7_16_r1 <= din_7_16;
    din_7_16_r2 <= din_7_16_r1;
    din_valid_7_17 <= out_new_pkt | hash_out_valid_filter_7_17;
    din_valid_7_17_r1 <= din_valid_7_17;
    din_valid_7_17_r2 <= din_valid_7_17_r1;

    din_7_17.data <= hash_out_valid_filter_7_17 ? hash_out_7_17 : 0;
    din_7_17.last <= out_new_pkt;
    din_7_17.bucket <= 7;


    din_7_17_r1 <= din_7_17;
    din_7_17_r2 <= din_7_17_r1;
    din_valid_7_18 <= out_new_pkt | hash_out_valid_filter_7_18;
    din_valid_7_18_r1 <= din_valid_7_18;
    din_valid_7_18_r2 <= din_valid_7_18_r1;

    din_7_18.data <= hash_out_valid_filter_7_18 ? hash_out_7_18 : 0;
    din_7_18.last <= out_new_pkt;
    din_7_18.bucket <= 7;


    din_7_18_r1 <= din_7_18;
    din_7_18_r2 <= din_7_18_r1;
    din_valid_7_19 <= out_new_pkt | hash_out_valid_filter_7_19;
    din_valid_7_19_r1 <= din_valid_7_19;
    din_valid_7_19_r2 <= din_valid_7_19_r1;

    din_7_19.data <= hash_out_valid_filter_7_19 ? hash_out_7_19 : 0;
    din_7_19.last <= out_new_pkt;
    din_7_19.bucket <= 7;


    din_7_19_r1 <= din_7_19;
    din_7_19_r2 <= din_7_19_r1;
    din_valid_7_20 <= out_new_pkt | hash_out_valid_filter_7_20;
    din_valid_7_20_r1 <= din_valid_7_20;
    din_valid_7_20_r2 <= din_valid_7_20_r1;

    din_7_20.data <= hash_out_valid_filter_7_20 ? hash_out_7_20 : 0;
    din_7_20.last <= out_new_pkt;
    din_7_20.bucket <= 7;


    din_7_20_r1 <= din_7_20;
    din_7_20_r2 <= din_7_20_r1;
    din_valid_7_21 <= out_new_pkt | hash_out_valid_filter_7_21;
    din_valid_7_21_r1 <= din_valid_7_21;
    din_valid_7_21_r2 <= din_valid_7_21_r1;

    din_7_21.data <= hash_out_valid_filter_7_21 ? hash_out_7_21 : 0;
    din_7_21.last <= out_new_pkt;
    din_7_21.bucket <= 7;


    din_7_21_r1 <= din_7_21;
    din_7_21_r2 <= din_7_21_r1;
    din_valid_7_22 <= out_new_pkt | hash_out_valid_filter_7_22;
    din_valid_7_22_r1 <= din_valid_7_22;
    din_valid_7_22_r2 <= din_valid_7_22_r1;

    din_7_22.data <= hash_out_valid_filter_7_22 ? hash_out_7_22 : 0;
    din_7_22.last <= out_new_pkt;
    din_7_22.bucket <= 7;


    din_7_22_r1 <= din_7_22;
    din_7_22_r2 <= din_7_22_r1;
    din_valid_7_23 <= out_new_pkt | hash_out_valid_filter_7_23;
    din_valid_7_23_r1 <= din_valid_7_23;
    din_valid_7_23_r2 <= din_valid_7_23_r1;

    din_7_23.data <= hash_out_valid_filter_7_23 ? hash_out_7_23 : 0;
    din_7_23.last <= out_new_pkt;
    din_7_23.bucket <= 7;


    din_7_23_r1 <= din_7_23;
    din_7_23_r2 <= din_7_23_r1;
    din_valid_7_24 <= out_new_pkt | hash_out_valid_filter_7_24;
    din_valid_7_24_r1 <= din_valid_7_24;
    din_valid_7_24_r2 <= din_valid_7_24_r1;

    din_7_24.data <= hash_out_valid_filter_7_24 ? hash_out_7_24 : 0;
    din_7_24.last <= out_new_pkt;
    din_7_24.bucket <= 7;


    din_7_24_r1 <= din_7_24;
    din_7_24_r2 <= din_7_24_r1;
    din_valid_7_25 <= out_new_pkt | hash_out_valid_filter_7_25;
    din_valid_7_25_r1 <= din_valid_7_25;
    din_valid_7_25_r2 <= din_valid_7_25_r1;

    din_7_25.data <= hash_out_valid_filter_7_25 ? hash_out_7_25 : 0;
    din_7_25.last <= out_new_pkt;
    din_7_25.bucket <= 7;


    din_7_25_r1 <= din_7_25;
    din_7_25_r2 <= din_7_25_r1;
    din_valid_7_26 <= out_new_pkt | hash_out_valid_filter_7_26;
    din_valid_7_26_r1 <= din_valid_7_26;
    din_valid_7_26_r2 <= din_valid_7_26_r1;

    din_7_26.data <= hash_out_valid_filter_7_26 ? hash_out_7_26 : 0;
    din_7_26.last <= out_new_pkt;
    din_7_26.bucket <= 7;


    din_7_26_r1 <= din_7_26;
    din_7_26_r2 <= din_7_26_r1;
    din_valid_7_27 <= out_new_pkt | hash_out_valid_filter_7_27;
    din_valid_7_27_r1 <= din_valid_7_27;
    din_valid_7_27_r2 <= din_valid_7_27_r1;

    din_7_27.data <= hash_out_valid_filter_7_27 ? hash_out_7_27 : 0;
    din_7_27.last <= out_new_pkt;
    din_7_27.bucket <= 7;


    din_7_27_r1 <= din_7_27;
    din_7_27_r2 <= din_7_27_r1;
    din_valid_7_28 <= out_new_pkt | hash_out_valid_filter_7_28;
    din_valid_7_28_r1 <= din_valid_7_28;
    din_valid_7_28_r2 <= din_valid_7_28_r1;

    din_7_28.data <= hash_out_valid_filter_7_28 ? hash_out_7_28 : 0;
    din_7_28.last <= out_new_pkt;
    din_7_28.bucket <= 7;


    din_7_28_r1 <= din_7_28;
    din_7_28_r2 <= din_7_28_r1;
    din_valid_7_29 <= out_new_pkt | hash_out_valid_filter_7_29;
    din_valid_7_29_r1 <= din_valid_7_29;
    din_valid_7_29_r2 <= din_valid_7_29_r1;

    din_7_29.data <= hash_out_valid_filter_7_29 ? hash_out_7_29 : 0;
    din_7_29.last <= out_new_pkt;
    din_7_29.bucket <= 7;


    din_7_29_r1 <= din_7_29;
    din_7_29_r2 <= din_7_29_r1;
    din_valid_7_30 <= out_new_pkt | hash_out_valid_filter_7_30;
    din_valid_7_30_r1 <= din_valid_7_30;
    din_valid_7_30_r2 <= din_valid_7_30_r1;

    din_7_30.data <= hash_out_valid_filter_7_30 ? hash_out_7_30 : 0;
    din_7_30.last <= out_new_pkt;
    din_7_30.bucket <= 7;


    din_7_30_r1 <= din_7_30;
    din_7_30_r2 <= din_7_30_r1;
    din_valid_7_31 <= out_new_pkt | hash_out_valid_filter_7_31;
    din_valid_7_31_r1 <= din_valid_7_31;
    din_valid_7_31_r2 <= din_valid_7_31_r1;

    din_7_31.data <= hash_out_valid_filter_7_31 ? hash_out_7_31 : 0;
    din_7_31.last <= out_new_pkt;
    din_7_31.bucket <= 7;


    din_7_31_r1 <= din_7_31;
    din_7_31_r2 <= din_7_31_r1;
end

//Instantiation
pkt_almost_full #(
    .DWIDTH(FP_DWIDTH),
    .EWIDTH(FP_EWIDTH),
    .NUM_PIPES(2)
) pkt_almost_full_inst (
    .clk                    (front_clk),
    .rst                    (front_rst),
    .in_data                (in_pkt_data),
    .in_valid               (in_pkt_valid),
    .in_ready               (in_pkt_ready),
    .in_sop                 (in_pkt_sop),
    .in_eop                 (in_pkt_eop),
    .in_empty               (in_pkt_empty),
    .out_data               (piped_pkt_data),
    .out_valid              (piped_pkt_valid),
    //.out_ready              (piped_pkt_ready),
    .out_almost_full        (piped_pkt_almost_full),
    .out_sop                (piped_pkt_sop),
    .out_eop                (piped_pkt_eop),
    .out_empty              (piped_pkt_empty)
);


frontend front(
    .clk(front_clk),
    .rst(front_rst),
    .hash_out_0_0 (hash_out_0_0),
    .hash_out_valid_filter_0_0(hash_out_valid_filter_0_0),
    .hash_out_0_1 (hash_out_0_1),
    .hash_out_valid_filter_0_1(hash_out_valid_filter_0_1),
    .hash_out_0_2 (hash_out_0_2),
    .hash_out_valid_filter_0_2(hash_out_valid_filter_0_2),
    .hash_out_0_3 (hash_out_0_3),
    .hash_out_valid_filter_0_3(hash_out_valid_filter_0_3),
    .hash_out_0_4 (hash_out_0_4),
    .hash_out_valid_filter_0_4(hash_out_valid_filter_0_4),
    .hash_out_0_5 (hash_out_0_5),
    .hash_out_valid_filter_0_5(hash_out_valid_filter_0_5),
    .hash_out_0_6 (hash_out_0_6),
    .hash_out_valid_filter_0_6(hash_out_valid_filter_0_6),
    .hash_out_0_7 (hash_out_0_7),
    .hash_out_valid_filter_0_7(hash_out_valid_filter_0_7),
    .hash_out_0_8 (hash_out_0_8),
    .hash_out_valid_filter_0_8(hash_out_valid_filter_0_8),
    .hash_out_0_9 (hash_out_0_9),
    .hash_out_valid_filter_0_9(hash_out_valid_filter_0_9),
    .hash_out_0_10 (hash_out_0_10),
    .hash_out_valid_filter_0_10(hash_out_valid_filter_0_10),
    .hash_out_0_11 (hash_out_0_11),
    .hash_out_valid_filter_0_11(hash_out_valid_filter_0_11),
    .hash_out_0_12 (hash_out_0_12),
    .hash_out_valid_filter_0_12(hash_out_valid_filter_0_12),
    .hash_out_0_13 (hash_out_0_13),
    .hash_out_valid_filter_0_13(hash_out_valid_filter_0_13),
    .hash_out_0_14 (hash_out_0_14),
    .hash_out_valid_filter_0_14(hash_out_valid_filter_0_14),
    .hash_out_0_15 (hash_out_0_15),
    .hash_out_valid_filter_0_15(hash_out_valid_filter_0_15),
    .hash_out_0_16 (hash_out_0_16),
    .hash_out_valid_filter_0_16(hash_out_valid_filter_0_16),
    .hash_out_0_17 (hash_out_0_17),
    .hash_out_valid_filter_0_17(hash_out_valid_filter_0_17),
    .hash_out_0_18 (hash_out_0_18),
    .hash_out_valid_filter_0_18(hash_out_valid_filter_0_18),
    .hash_out_0_19 (hash_out_0_19),
    .hash_out_valid_filter_0_19(hash_out_valid_filter_0_19),
    .hash_out_0_20 (hash_out_0_20),
    .hash_out_valid_filter_0_20(hash_out_valid_filter_0_20),
    .hash_out_0_21 (hash_out_0_21),
    .hash_out_valid_filter_0_21(hash_out_valid_filter_0_21),
    .hash_out_0_22 (hash_out_0_22),
    .hash_out_valid_filter_0_22(hash_out_valid_filter_0_22),
    .hash_out_0_23 (hash_out_0_23),
    .hash_out_valid_filter_0_23(hash_out_valid_filter_0_23),
    .hash_out_0_24 (hash_out_0_24),
    .hash_out_valid_filter_0_24(hash_out_valid_filter_0_24),
    .hash_out_0_25 (hash_out_0_25),
    .hash_out_valid_filter_0_25(hash_out_valid_filter_0_25),
    .hash_out_0_26 (hash_out_0_26),
    .hash_out_valid_filter_0_26(hash_out_valid_filter_0_26),
    .hash_out_0_27 (hash_out_0_27),
    .hash_out_valid_filter_0_27(hash_out_valid_filter_0_27),
    .hash_out_0_28 (hash_out_0_28),
    .hash_out_valid_filter_0_28(hash_out_valid_filter_0_28),
    .hash_out_0_29 (hash_out_0_29),
    .hash_out_valid_filter_0_29(hash_out_valid_filter_0_29),
    .hash_out_0_30 (hash_out_0_30),
    .hash_out_valid_filter_0_30(hash_out_valid_filter_0_30),
    .hash_out_0_31 (hash_out_0_31),
    .hash_out_valid_filter_0_31(hash_out_valid_filter_0_31),
    .hash_out_1_0 (hash_out_1_0),
    .hash_out_valid_filter_1_0(hash_out_valid_filter_1_0),
    .hash_out_1_1 (hash_out_1_1),
    .hash_out_valid_filter_1_1(hash_out_valid_filter_1_1),
    .hash_out_1_2 (hash_out_1_2),
    .hash_out_valid_filter_1_2(hash_out_valid_filter_1_2),
    .hash_out_1_3 (hash_out_1_3),
    .hash_out_valid_filter_1_3(hash_out_valid_filter_1_3),
    .hash_out_1_4 (hash_out_1_4),
    .hash_out_valid_filter_1_4(hash_out_valid_filter_1_4),
    .hash_out_1_5 (hash_out_1_5),
    .hash_out_valid_filter_1_5(hash_out_valid_filter_1_5),
    .hash_out_1_6 (hash_out_1_6),
    .hash_out_valid_filter_1_6(hash_out_valid_filter_1_6),
    .hash_out_1_7 (hash_out_1_7),
    .hash_out_valid_filter_1_7(hash_out_valid_filter_1_7),
    .hash_out_1_8 (hash_out_1_8),
    .hash_out_valid_filter_1_8(hash_out_valid_filter_1_8),
    .hash_out_1_9 (hash_out_1_9),
    .hash_out_valid_filter_1_9(hash_out_valid_filter_1_9),
    .hash_out_1_10 (hash_out_1_10),
    .hash_out_valid_filter_1_10(hash_out_valid_filter_1_10),
    .hash_out_1_11 (hash_out_1_11),
    .hash_out_valid_filter_1_11(hash_out_valid_filter_1_11),
    .hash_out_1_12 (hash_out_1_12),
    .hash_out_valid_filter_1_12(hash_out_valid_filter_1_12),
    .hash_out_1_13 (hash_out_1_13),
    .hash_out_valid_filter_1_13(hash_out_valid_filter_1_13),
    .hash_out_1_14 (hash_out_1_14),
    .hash_out_valid_filter_1_14(hash_out_valid_filter_1_14),
    .hash_out_1_15 (hash_out_1_15),
    .hash_out_valid_filter_1_15(hash_out_valid_filter_1_15),
    .hash_out_1_16 (hash_out_1_16),
    .hash_out_valid_filter_1_16(hash_out_valid_filter_1_16),
    .hash_out_1_17 (hash_out_1_17),
    .hash_out_valid_filter_1_17(hash_out_valid_filter_1_17),
    .hash_out_1_18 (hash_out_1_18),
    .hash_out_valid_filter_1_18(hash_out_valid_filter_1_18),
    .hash_out_1_19 (hash_out_1_19),
    .hash_out_valid_filter_1_19(hash_out_valid_filter_1_19),
    .hash_out_1_20 (hash_out_1_20),
    .hash_out_valid_filter_1_20(hash_out_valid_filter_1_20),
    .hash_out_1_21 (hash_out_1_21),
    .hash_out_valid_filter_1_21(hash_out_valid_filter_1_21),
    .hash_out_1_22 (hash_out_1_22),
    .hash_out_valid_filter_1_22(hash_out_valid_filter_1_22),
    .hash_out_1_23 (hash_out_1_23),
    .hash_out_valid_filter_1_23(hash_out_valid_filter_1_23),
    .hash_out_1_24 (hash_out_1_24),
    .hash_out_valid_filter_1_24(hash_out_valid_filter_1_24),
    .hash_out_1_25 (hash_out_1_25),
    .hash_out_valid_filter_1_25(hash_out_valid_filter_1_25),
    .hash_out_1_26 (hash_out_1_26),
    .hash_out_valid_filter_1_26(hash_out_valid_filter_1_26),
    .hash_out_1_27 (hash_out_1_27),
    .hash_out_valid_filter_1_27(hash_out_valid_filter_1_27),
    .hash_out_1_28 (hash_out_1_28),
    .hash_out_valid_filter_1_28(hash_out_valid_filter_1_28),
    .hash_out_1_29 (hash_out_1_29),
    .hash_out_valid_filter_1_29(hash_out_valid_filter_1_29),
    .hash_out_1_30 (hash_out_1_30),
    .hash_out_valid_filter_1_30(hash_out_valid_filter_1_30),
    .hash_out_1_31 (hash_out_1_31),
    .hash_out_valid_filter_1_31(hash_out_valid_filter_1_31),
    .hash_out_2_0 (hash_out_2_0),
    .hash_out_valid_filter_2_0(hash_out_valid_filter_2_0),
    .hash_out_2_1 (hash_out_2_1),
    .hash_out_valid_filter_2_1(hash_out_valid_filter_2_1),
    .hash_out_2_2 (hash_out_2_2),
    .hash_out_valid_filter_2_2(hash_out_valid_filter_2_2),
    .hash_out_2_3 (hash_out_2_3),
    .hash_out_valid_filter_2_3(hash_out_valid_filter_2_3),
    .hash_out_2_4 (hash_out_2_4),
    .hash_out_valid_filter_2_4(hash_out_valid_filter_2_4),
    .hash_out_2_5 (hash_out_2_5),
    .hash_out_valid_filter_2_5(hash_out_valid_filter_2_5),
    .hash_out_2_6 (hash_out_2_6),
    .hash_out_valid_filter_2_6(hash_out_valid_filter_2_6),
    .hash_out_2_7 (hash_out_2_7),
    .hash_out_valid_filter_2_7(hash_out_valid_filter_2_7),
    .hash_out_2_8 (hash_out_2_8),
    .hash_out_valid_filter_2_8(hash_out_valid_filter_2_8),
    .hash_out_2_9 (hash_out_2_9),
    .hash_out_valid_filter_2_9(hash_out_valid_filter_2_9),
    .hash_out_2_10 (hash_out_2_10),
    .hash_out_valid_filter_2_10(hash_out_valid_filter_2_10),
    .hash_out_2_11 (hash_out_2_11),
    .hash_out_valid_filter_2_11(hash_out_valid_filter_2_11),
    .hash_out_2_12 (hash_out_2_12),
    .hash_out_valid_filter_2_12(hash_out_valid_filter_2_12),
    .hash_out_2_13 (hash_out_2_13),
    .hash_out_valid_filter_2_13(hash_out_valid_filter_2_13),
    .hash_out_2_14 (hash_out_2_14),
    .hash_out_valid_filter_2_14(hash_out_valid_filter_2_14),
    .hash_out_2_15 (hash_out_2_15),
    .hash_out_valid_filter_2_15(hash_out_valid_filter_2_15),
    .hash_out_2_16 (hash_out_2_16),
    .hash_out_valid_filter_2_16(hash_out_valid_filter_2_16),
    .hash_out_2_17 (hash_out_2_17),
    .hash_out_valid_filter_2_17(hash_out_valid_filter_2_17),
    .hash_out_2_18 (hash_out_2_18),
    .hash_out_valid_filter_2_18(hash_out_valid_filter_2_18),
    .hash_out_2_19 (hash_out_2_19),
    .hash_out_valid_filter_2_19(hash_out_valid_filter_2_19),
    .hash_out_2_20 (hash_out_2_20),
    .hash_out_valid_filter_2_20(hash_out_valid_filter_2_20),
    .hash_out_2_21 (hash_out_2_21),
    .hash_out_valid_filter_2_21(hash_out_valid_filter_2_21),
    .hash_out_2_22 (hash_out_2_22),
    .hash_out_valid_filter_2_22(hash_out_valid_filter_2_22),
    .hash_out_2_23 (hash_out_2_23),
    .hash_out_valid_filter_2_23(hash_out_valid_filter_2_23),
    .hash_out_2_24 (hash_out_2_24),
    .hash_out_valid_filter_2_24(hash_out_valid_filter_2_24),
    .hash_out_2_25 (hash_out_2_25),
    .hash_out_valid_filter_2_25(hash_out_valid_filter_2_25),
    .hash_out_2_26 (hash_out_2_26),
    .hash_out_valid_filter_2_26(hash_out_valid_filter_2_26),
    .hash_out_2_27 (hash_out_2_27),
    .hash_out_valid_filter_2_27(hash_out_valid_filter_2_27),
    .hash_out_2_28 (hash_out_2_28),
    .hash_out_valid_filter_2_28(hash_out_valid_filter_2_28),
    .hash_out_2_29 (hash_out_2_29),
    .hash_out_valid_filter_2_29(hash_out_valid_filter_2_29),
    .hash_out_2_30 (hash_out_2_30),
    .hash_out_valid_filter_2_30(hash_out_valid_filter_2_30),
    .hash_out_2_31 (hash_out_2_31),
    .hash_out_valid_filter_2_31(hash_out_valid_filter_2_31),
    .hash_out_3_0 (hash_out_3_0),
    .hash_out_valid_filter_3_0(hash_out_valid_filter_3_0),
    .hash_out_3_1 (hash_out_3_1),
    .hash_out_valid_filter_3_1(hash_out_valid_filter_3_1),
    .hash_out_3_2 (hash_out_3_2),
    .hash_out_valid_filter_3_2(hash_out_valid_filter_3_2),
    .hash_out_3_3 (hash_out_3_3),
    .hash_out_valid_filter_3_3(hash_out_valid_filter_3_3),
    .hash_out_3_4 (hash_out_3_4),
    .hash_out_valid_filter_3_4(hash_out_valid_filter_3_4),
    .hash_out_3_5 (hash_out_3_5),
    .hash_out_valid_filter_3_5(hash_out_valid_filter_3_5),
    .hash_out_3_6 (hash_out_3_6),
    .hash_out_valid_filter_3_6(hash_out_valid_filter_3_6),
    .hash_out_3_7 (hash_out_3_7),
    .hash_out_valid_filter_3_7(hash_out_valid_filter_3_7),
    .hash_out_3_8 (hash_out_3_8),
    .hash_out_valid_filter_3_8(hash_out_valid_filter_3_8),
    .hash_out_3_9 (hash_out_3_9),
    .hash_out_valid_filter_3_9(hash_out_valid_filter_3_9),
    .hash_out_3_10 (hash_out_3_10),
    .hash_out_valid_filter_3_10(hash_out_valid_filter_3_10),
    .hash_out_3_11 (hash_out_3_11),
    .hash_out_valid_filter_3_11(hash_out_valid_filter_3_11),
    .hash_out_3_12 (hash_out_3_12),
    .hash_out_valid_filter_3_12(hash_out_valid_filter_3_12),
    .hash_out_3_13 (hash_out_3_13),
    .hash_out_valid_filter_3_13(hash_out_valid_filter_3_13),
    .hash_out_3_14 (hash_out_3_14),
    .hash_out_valid_filter_3_14(hash_out_valid_filter_3_14),
    .hash_out_3_15 (hash_out_3_15),
    .hash_out_valid_filter_3_15(hash_out_valid_filter_3_15),
    .hash_out_3_16 (hash_out_3_16),
    .hash_out_valid_filter_3_16(hash_out_valid_filter_3_16),
    .hash_out_3_17 (hash_out_3_17),
    .hash_out_valid_filter_3_17(hash_out_valid_filter_3_17),
    .hash_out_3_18 (hash_out_3_18),
    .hash_out_valid_filter_3_18(hash_out_valid_filter_3_18),
    .hash_out_3_19 (hash_out_3_19),
    .hash_out_valid_filter_3_19(hash_out_valid_filter_3_19),
    .hash_out_3_20 (hash_out_3_20),
    .hash_out_valid_filter_3_20(hash_out_valid_filter_3_20),
    .hash_out_3_21 (hash_out_3_21),
    .hash_out_valid_filter_3_21(hash_out_valid_filter_3_21),
    .hash_out_3_22 (hash_out_3_22),
    .hash_out_valid_filter_3_22(hash_out_valid_filter_3_22),
    .hash_out_3_23 (hash_out_3_23),
    .hash_out_valid_filter_3_23(hash_out_valid_filter_3_23),
    .hash_out_3_24 (hash_out_3_24),
    .hash_out_valid_filter_3_24(hash_out_valid_filter_3_24),
    .hash_out_3_25 (hash_out_3_25),
    .hash_out_valid_filter_3_25(hash_out_valid_filter_3_25),
    .hash_out_3_26 (hash_out_3_26),
    .hash_out_valid_filter_3_26(hash_out_valid_filter_3_26),
    .hash_out_3_27 (hash_out_3_27),
    .hash_out_valid_filter_3_27(hash_out_valid_filter_3_27),
    .hash_out_3_28 (hash_out_3_28),
    .hash_out_valid_filter_3_28(hash_out_valid_filter_3_28),
    .hash_out_3_29 (hash_out_3_29),
    .hash_out_valid_filter_3_29(hash_out_valid_filter_3_29),
    .hash_out_3_30 (hash_out_3_30),
    .hash_out_valid_filter_3_30(hash_out_valid_filter_3_30),
    .hash_out_3_31 (hash_out_3_31),
    .hash_out_valid_filter_3_31(hash_out_valid_filter_3_31),
    .hash_out_4_0 (hash_out_4_0),
    .hash_out_valid_filter_4_0(hash_out_valid_filter_4_0),
    .hash_out_4_1 (hash_out_4_1),
    .hash_out_valid_filter_4_1(hash_out_valid_filter_4_1),
    .hash_out_4_2 (hash_out_4_2),
    .hash_out_valid_filter_4_2(hash_out_valid_filter_4_2),
    .hash_out_4_3 (hash_out_4_3),
    .hash_out_valid_filter_4_3(hash_out_valid_filter_4_3),
    .hash_out_4_4 (hash_out_4_4),
    .hash_out_valid_filter_4_4(hash_out_valid_filter_4_4),
    .hash_out_4_5 (hash_out_4_5),
    .hash_out_valid_filter_4_5(hash_out_valid_filter_4_5),
    .hash_out_4_6 (hash_out_4_6),
    .hash_out_valid_filter_4_6(hash_out_valid_filter_4_6),
    .hash_out_4_7 (hash_out_4_7),
    .hash_out_valid_filter_4_7(hash_out_valid_filter_4_7),
    .hash_out_4_8 (hash_out_4_8),
    .hash_out_valid_filter_4_8(hash_out_valid_filter_4_8),
    .hash_out_4_9 (hash_out_4_9),
    .hash_out_valid_filter_4_9(hash_out_valid_filter_4_9),
    .hash_out_4_10 (hash_out_4_10),
    .hash_out_valid_filter_4_10(hash_out_valid_filter_4_10),
    .hash_out_4_11 (hash_out_4_11),
    .hash_out_valid_filter_4_11(hash_out_valid_filter_4_11),
    .hash_out_4_12 (hash_out_4_12),
    .hash_out_valid_filter_4_12(hash_out_valid_filter_4_12),
    .hash_out_4_13 (hash_out_4_13),
    .hash_out_valid_filter_4_13(hash_out_valid_filter_4_13),
    .hash_out_4_14 (hash_out_4_14),
    .hash_out_valid_filter_4_14(hash_out_valid_filter_4_14),
    .hash_out_4_15 (hash_out_4_15),
    .hash_out_valid_filter_4_15(hash_out_valid_filter_4_15),
    .hash_out_4_16 (hash_out_4_16),
    .hash_out_valid_filter_4_16(hash_out_valid_filter_4_16),
    .hash_out_4_17 (hash_out_4_17),
    .hash_out_valid_filter_4_17(hash_out_valid_filter_4_17),
    .hash_out_4_18 (hash_out_4_18),
    .hash_out_valid_filter_4_18(hash_out_valid_filter_4_18),
    .hash_out_4_19 (hash_out_4_19),
    .hash_out_valid_filter_4_19(hash_out_valid_filter_4_19),
    .hash_out_4_20 (hash_out_4_20),
    .hash_out_valid_filter_4_20(hash_out_valid_filter_4_20),
    .hash_out_4_21 (hash_out_4_21),
    .hash_out_valid_filter_4_21(hash_out_valid_filter_4_21),
    .hash_out_4_22 (hash_out_4_22),
    .hash_out_valid_filter_4_22(hash_out_valid_filter_4_22),
    .hash_out_4_23 (hash_out_4_23),
    .hash_out_valid_filter_4_23(hash_out_valid_filter_4_23),
    .hash_out_4_24 (hash_out_4_24),
    .hash_out_valid_filter_4_24(hash_out_valid_filter_4_24),
    .hash_out_4_25 (hash_out_4_25),
    .hash_out_valid_filter_4_25(hash_out_valid_filter_4_25),
    .hash_out_4_26 (hash_out_4_26),
    .hash_out_valid_filter_4_26(hash_out_valid_filter_4_26),
    .hash_out_4_27 (hash_out_4_27),
    .hash_out_valid_filter_4_27(hash_out_valid_filter_4_27),
    .hash_out_4_28 (hash_out_4_28),
    .hash_out_valid_filter_4_28(hash_out_valid_filter_4_28),
    .hash_out_4_29 (hash_out_4_29),
    .hash_out_valid_filter_4_29(hash_out_valid_filter_4_29),
    .hash_out_4_30 (hash_out_4_30),
    .hash_out_valid_filter_4_30(hash_out_valid_filter_4_30),
    .hash_out_4_31 (hash_out_4_31),
    .hash_out_valid_filter_4_31(hash_out_valid_filter_4_31),
    .hash_out_5_0 (hash_out_5_0),
    .hash_out_valid_filter_5_0(hash_out_valid_filter_5_0),
    .hash_out_5_1 (hash_out_5_1),
    .hash_out_valid_filter_5_1(hash_out_valid_filter_5_1),
    .hash_out_5_2 (hash_out_5_2),
    .hash_out_valid_filter_5_2(hash_out_valid_filter_5_2),
    .hash_out_5_3 (hash_out_5_3),
    .hash_out_valid_filter_5_3(hash_out_valid_filter_5_3),
    .hash_out_5_4 (hash_out_5_4),
    .hash_out_valid_filter_5_4(hash_out_valid_filter_5_4),
    .hash_out_5_5 (hash_out_5_5),
    .hash_out_valid_filter_5_5(hash_out_valid_filter_5_5),
    .hash_out_5_6 (hash_out_5_6),
    .hash_out_valid_filter_5_6(hash_out_valid_filter_5_6),
    .hash_out_5_7 (hash_out_5_7),
    .hash_out_valid_filter_5_7(hash_out_valid_filter_5_7),
    .hash_out_5_8 (hash_out_5_8),
    .hash_out_valid_filter_5_8(hash_out_valid_filter_5_8),
    .hash_out_5_9 (hash_out_5_9),
    .hash_out_valid_filter_5_9(hash_out_valid_filter_5_9),
    .hash_out_5_10 (hash_out_5_10),
    .hash_out_valid_filter_5_10(hash_out_valid_filter_5_10),
    .hash_out_5_11 (hash_out_5_11),
    .hash_out_valid_filter_5_11(hash_out_valid_filter_5_11),
    .hash_out_5_12 (hash_out_5_12),
    .hash_out_valid_filter_5_12(hash_out_valid_filter_5_12),
    .hash_out_5_13 (hash_out_5_13),
    .hash_out_valid_filter_5_13(hash_out_valid_filter_5_13),
    .hash_out_5_14 (hash_out_5_14),
    .hash_out_valid_filter_5_14(hash_out_valid_filter_5_14),
    .hash_out_5_15 (hash_out_5_15),
    .hash_out_valid_filter_5_15(hash_out_valid_filter_5_15),
    .hash_out_5_16 (hash_out_5_16),
    .hash_out_valid_filter_5_16(hash_out_valid_filter_5_16),
    .hash_out_5_17 (hash_out_5_17),
    .hash_out_valid_filter_5_17(hash_out_valid_filter_5_17),
    .hash_out_5_18 (hash_out_5_18),
    .hash_out_valid_filter_5_18(hash_out_valid_filter_5_18),
    .hash_out_5_19 (hash_out_5_19),
    .hash_out_valid_filter_5_19(hash_out_valid_filter_5_19),
    .hash_out_5_20 (hash_out_5_20),
    .hash_out_valid_filter_5_20(hash_out_valid_filter_5_20),
    .hash_out_5_21 (hash_out_5_21),
    .hash_out_valid_filter_5_21(hash_out_valid_filter_5_21),
    .hash_out_5_22 (hash_out_5_22),
    .hash_out_valid_filter_5_22(hash_out_valid_filter_5_22),
    .hash_out_5_23 (hash_out_5_23),
    .hash_out_valid_filter_5_23(hash_out_valid_filter_5_23),
    .hash_out_5_24 (hash_out_5_24),
    .hash_out_valid_filter_5_24(hash_out_valid_filter_5_24),
    .hash_out_5_25 (hash_out_5_25),
    .hash_out_valid_filter_5_25(hash_out_valid_filter_5_25),
    .hash_out_5_26 (hash_out_5_26),
    .hash_out_valid_filter_5_26(hash_out_valid_filter_5_26),
    .hash_out_5_27 (hash_out_5_27),
    .hash_out_valid_filter_5_27(hash_out_valid_filter_5_27),
    .hash_out_5_28 (hash_out_5_28),
    .hash_out_valid_filter_5_28(hash_out_valid_filter_5_28),
    .hash_out_5_29 (hash_out_5_29),
    .hash_out_valid_filter_5_29(hash_out_valid_filter_5_29),
    .hash_out_5_30 (hash_out_5_30),
    .hash_out_valid_filter_5_30(hash_out_valid_filter_5_30),
    .hash_out_5_31 (hash_out_5_31),
    .hash_out_valid_filter_5_31(hash_out_valid_filter_5_31),
    .hash_out_6_0 (hash_out_6_0),
    .hash_out_valid_filter_6_0(hash_out_valid_filter_6_0),
    .hash_out_6_1 (hash_out_6_1),
    .hash_out_valid_filter_6_1(hash_out_valid_filter_6_1),
    .hash_out_6_2 (hash_out_6_2),
    .hash_out_valid_filter_6_2(hash_out_valid_filter_6_2),
    .hash_out_6_3 (hash_out_6_3),
    .hash_out_valid_filter_6_3(hash_out_valid_filter_6_3),
    .hash_out_6_4 (hash_out_6_4),
    .hash_out_valid_filter_6_4(hash_out_valid_filter_6_4),
    .hash_out_6_5 (hash_out_6_5),
    .hash_out_valid_filter_6_5(hash_out_valid_filter_6_5),
    .hash_out_6_6 (hash_out_6_6),
    .hash_out_valid_filter_6_6(hash_out_valid_filter_6_6),
    .hash_out_6_7 (hash_out_6_7),
    .hash_out_valid_filter_6_7(hash_out_valid_filter_6_7),
    .hash_out_6_8 (hash_out_6_8),
    .hash_out_valid_filter_6_8(hash_out_valid_filter_6_8),
    .hash_out_6_9 (hash_out_6_9),
    .hash_out_valid_filter_6_9(hash_out_valid_filter_6_9),
    .hash_out_6_10 (hash_out_6_10),
    .hash_out_valid_filter_6_10(hash_out_valid_filter_6_10),
    .hash_out_6_11 (hash_out_6_11),
    .hash_out_valid_filter_6_11(hash_out_valid_filter_6_11),
    .hash_out_6_12 (hash_out_6_12),
    .hash_out_valid_filter_6_12(hash_out_valid_filter_6_12),
    .hash_out_6_13 (hash_out_6_13),
    .hash_out_valid_filter_6_13(hash_out_valid_filter_6_13),
    .hash_out_6_14 (hash_out_6_14),
    .hash_out_valid_filter_6_14(hash_out_valid_filter_6_14),
    .hash_out_6_15 (hash_out_6_15),
    .hash_out_valid_filter_6_15(hash_out_valid_filter_6_15),
    .hash_out_6_16 (hash_out_6_16),
    .hash_out_valid_filter_6_16(hash_out_valid_filter_6_16),
    .hash_out_6_17 (hash_out_6_17),
    .hash_out_valid_filter_6_17(hash_out_valid_filter_6_17),
    .hash_out_6_18 (hash_out_6_18),
    .hash_out_valid_filter_6_18(hash_out_valid_filter_6_18),
    .hash_out_6_19 (hash_out_6_19),
    .hash_out_valid_filter_6_19(hash_out_valid_filter_6_19),
    .hash_out_6_20 (hash_out_6_20),
    .hash_out_valid_filter_6_20(hash_out_valid_filter_6_20),
    .hash_out_6_21 (hash_out_6_21),
    .hash_out_valid_filter_6_21(hash_out_valid_filter_6_21),
    .hash_out_6_22 (hash_out_6_22),
    .hash_out_valid_filter_6_22(hash_out_valid_filter_6_22),
    .hash_out_6_23 (hash_out_6_23),
    .hash_out_valid_filter_6_23(hash_out_valid_filter_6_23),
    .hash_out_6_24 (hash_out_6_24),
    .hash_out_valid_filter_6_24(hash_out_valid_filter_6_24),
    .hash_out_6_25 (hash_out_6_25),
    .hash_out_valid_filter_6_25(hash_out_valid_filter_6_25),
    .hash_out_6_26 (hash_out_6_26),
    .hash_out_valid_filter_6_26(hash_out_valid_filter_6_26),
    .hash_out_6_27 (hash_out_6_27),
    .hash_out_valid_filter_6_27(hash_out_valid_filter_6_27),
    .hash_out_6_28 (hash_out_6_28),
    .hash_out_valid_filter_6_28(hash_out_valid_filter_6_28),
    .hash_out_6_29 (hash_out_6_29),
    .hash_out_valid_filter_6_29(hash_out_valid_filter_6_29),
    .hash_out_6_30 (hash_out_6_30),
    .hash_out_valid_filter_6_30(hash_out_valid_filter_6_30),
    .hash_out_6_31 (hash_out_6_31),
    .hash_out_valid_filter_6_31(hash_out_valid_filter_6_31),
    .hash_out_7_0 (hash_out_7_0),
    .hash_out_valid_filter_7_0(hash_out_valid_filter_7_0),
    .hash_out_7_1 (hash_out_7_1),
    .hash_out_valid_filter_7_1(hash_out_valid_filter_7_1),
    .hash_out_7_2 (hash_out_7_2),
    .hash_out_valid_filter_7_2(hash_out_valid_filter_7_2),
    .hash_out_7_3 (hash_out_7_3),
    .hash_out_valid_filter_7_3(hash_out_valid_filter_7_3),
    .hash_out_7_4 (hash_out_7_4),
    .hash_out_valid_filter_7_4(hash_out_valid_filter_7_4),
    .hash_out_7_5 (hash_out_7_5),
    .hash_out_valid_filter_7_5(hash_out_valid_filter_7_5),
    .hash_out_7_6 (hash_out_7_6),
    .hash_out_valid_filter_7_6(hash_out_valid_filter_7_6),
    .hash_out_7_7 (hash_out_7_7),
    .hash_out_valid_filter_7_7(hash_out_valid_filter_7_7),
    .hash_out_7_8 (hash_out_7_8),
    .hash_out_valid_filter_7_8(hash_out_valid_filter_7_8),
    .hash_out_7_9 (hash_out_7_9),
    .hash_out_valid_filter_7_9(hash_out_valid_filter_7_9),
    .hash_out_7_10 (hash_out_7_10),
    .hash_out_valid_filter_7_10(hash_out_valid_filter_7_10),
    .hash_out_7_11 (hash_out_7_11),
    .hash_out_valid_filter_7_11(hash_out_valid_filter_7_11),
    .hash_out_7_12 (hash_out_7_12),
    .hash_out_valid_filter_7_12(hash_out_valid_filter_7_12),
    .hash_out_7_13 (hash_out_7_13),
    .hash_out_valid_filter_7_13(hash_out_valid_filter_7_13),
    .hash_out_7_14 (hash_out_7_14),
    .hash_out_valid_filter_7_14(hash_out_valid_filter_7_14),
    .hash_out_7_15 (hash_out_7_15),
    .hash_out_valid_filter_7_15(hash_out_valid_filter_7_15),
    .hash_out_7_16 (hash_out_7_16),
    .hash_out_valid_filter_7_16(hash_out_valid_filter_7_16),
    .hash_out_7_17 (hash_out_7_17),
    .hash_out_valid_filter_7_17(hash_out_valid_filter_7_17),
    .hash_out_7_18 (hash_out_7_18),
    .hash_out_valid_filter_7_18(hash_out_valid_filter_7_18),
    .hash_out_7_19 (hash_out_7_19),
    .hash_out_valid_filter_7_19(hash_out_valid_filter_7_19),
    .hash_out_7_20 (hash_out_7_20),
    .hash_out_valid_filter_7_20(hash_out_valid_filter_7_20),
    .hash_out_7_21 (hash_out_7_21),
    .hash_out_valid_filter_7_21(hash_out_valid_filter_7_21),
    .hash_out_7_22 (hash_out_7_22),
    .hash_out_valid_filter_7_22(hash_out_valid_filter_7_22),
    .hash_out_7_23 (hash_out_7_23),
    .hash_out_valid_filter_7_23(hash_out_valid_filter_7_23),
    .hash_out_7_24 (hash_out_7_24),
    .hash_out_valid_filter_7_24(hash_out_valid_filter_7_24),
    .hash_out_7_25 (hash_out_7_25),
    .hash_out_valid_filter_7_25(hash_out_valid_filter_7_25),
    .hash_out_7_26 (hash_out_7_26),
    .hash_out_valid_filter_7_26(hash_out_valid_filter_7_26),
    .hash_out_7_27 (hash_out_7_27),
    .hash_out_valid_filter_7_27(hash_out_valid_filter_7_27),
    .hash_out_7_28 (hash_out_7_28),
    .hash_out_valid_filter_7_28(hash_out_valid_filter_7_28),
    .hash_out_7_29 (hash_out_7_29),
    .hash_out_valid_filter_7_29(hash_out_valid_filter_7_29),
    .hash_out_7_30 (hash_out_7_30),
    .hash_out_valid_filter_7_30(hash_out_valid_filter_7_30),
    .hash_out_7_31 (hash_out_7_31),
    .hash_out_valid_filter_7_31(hash_out_valid_filter_7_31),
    .in_data         (piped_pkt_data_swap),
    .in_valid        (piped_pkt_valid),
    .in_sop          (piped_pkt_sop),
    .in_eop          (piped_pkt_eop),
    .in_empty        (piped_pkt_empty),
    .out_new_pkt     (out_new_pkt)
);
//RuleID reduction logic
backend back(
    .clk                     (back_clk),
    .rst                     (back_rst),
    .in_data_0_0     (back_data_0_0),
    .in_valid_0_0    (back_valid_0_0),
    .in_ready_0_0    (back_ready_0_0),
    .in_data_0_1     (back_data_0_1),
    .in_valid_0_1    (back_valid_0_1),
    .in_ready_0_1    (back_ready_0_1),
    .in_data_0_2     (back_data_0_2),
    .in_valid_0_2    (back_valid_0_2),
    .in_ready_0_2    (back_ready_0_2),
    .in_data_0_3     (back_data_0_3),
    .in_valid_0_3    (back_valid_0_3),
    .in_ready_0_3    (back_ready_0_3),
    .in_data_0_4     (back_data_0_4),
    .in_valid_0_4    (back_valid_0_4),
    .in_ready_0_4    (back_ready_0_4),
    .in_data_0_5     (back_data_0_5),
    .in_valid_0_5    (back_valid_0_5),
    .in_ready_0_5    (back_ready_0_5),
    .in_data_0_6     (back_data_0_6),
    .in_valid_0_6    (back_valid_0_6),
    .in_ready_0_6    (back_ready_0_6),
    .in_data_0_7     (back_data_0_7),
    .in_valid_0_7    (back_valid_0_7),
    .in_ready_0_7    (back_ready_0_7),
    .in_data_0_8     (back_data_0_8),
    .in_valid_0_8    (back_valid_0_8),
    .in_ready_0_8    (back_ready_0_8),
    .in_data_0_9     (back_data_0_9),
    .in_valid_0_9    (back_valid_0_9),
    .in_ready_0_9    (back_ready_0_9),
    .in_data_0_10     (back_data_0_10),
    .in_valid_0_10    (back_valid_0_10),
    .in_ready_0_10    (back_ready_0_10),
    .in_data_0_11     (back_data_0_11),
    .in_valid_0_11    (back_valid_0_11),
    .in_ready_0_11    (back_ready_0_11),
    .in_data_0_12     (back_data_0_12),
    .in_valid_0_12    (back_valid_0_12),
    .in_ready_0_12    (back_ready_0_12),
    .in_data_0_13     (back_data_0_13),
    .in_valid_0_13    (back_valid_0_13),
    .in_ready_0_13    (back_ready_0_13),
    .in_data_0_14     (back_data_0_14),
    .in_valid_0_14    (back_valid_0_14),
    .in_ready_0_14    (back_ready_0_14),
    .in_data_0_15     (back_data_0_15),
    .in_valid_0_15    (back_valid_0_15),
    .in_ready_0_15    (back_ready_0_15),
    .in_data_0_16     (back_data_0_16),
    .in_valid_0_16    (back_valid_0_16),
    .in_ready_0_16    (back_ready_0_16),
    .in_data_0_17     (back_data_0_17),
    .in_valid_0_17    (back_valid_0_17),
    .in_ready_0_17    (back_ready_0_17),
    .in_data_0_18     (back_data_0_18),
    .in_valid_0_18    (back_valid_0_18),
    .in_ready_0_18    (back_ready_0_18),
    .in_data_0_19     (back_data_0_19),
    .in_valid_0_19    (back_valid_0_19),
    .in_ready_0_19    (back_ready_0_19),
    .in_data_0_20     (back_data_0_20),
    .in_valid_0_20    (back_valid_0_20),
    .in_ready_0_20    (back_ready_0_20),
    .in_data_0_21     (back_data_0_21),
    .in_valid_0_21    (back_valid_0_21),
    .in_ready_0_21    (back_ready_0_21),
    .in_data_0_22     (back_data_0_22),
    .in_valid_0_22    (back_valid_0_22),
    .in_ready_0_22    (back_ready_0_22),
    .in_data_0_23     (back_data_0_23),
    .in_valid_0_23    (back_valid_0_23),
    .in_ready_0_23    (back_ready_0_23),
    .in_data_0_24     (back_data_0_24),
    .in_valid_0_24    (back_valid_0_24),
    .in_ready_0_24    (back_ready_0_24),
    .in_data_0_25     (back_data_0_25),
    .in_valid_0_25    (back_valid_0_25),
    .in_ready_0_25    (back_ready_0_25),
    .in_data_0_26     (back_data_0_26),
    .in_valid_0_26    (back_valid_0_26),
    .in_ready_0_26    (back_ready_0_26),
    .in_data_0_27     (back_data_0_27),
    .in_valid_0_27    (back_valid_0_27),
    .in_ready_0_27    (back_ready_0_27),
    .in_data_0_28     (back_data_0_28),
    .in_valid_0_28    (back_valid_0_28),
    .in_ready_0_28    (back_ready_0_28),
    .in_data_0_29     (back_data_0_29),
    .in_valid_0_29    (back_valid_0_29),
    .in_ready_0_29    (back_ready_0_29),
    .in_data_0_30     (back_data_0_30),
    .in_valid_0_30    (back_valid_0_30),
    .in_ready_0_30    (back_ready_0_30),
    .in_data_0_31     (back_data_0_31),
    .in_valid_0_31    (back_valid_0_31),
    .in_ready_0_31    (back_ready_0_31),
    .in_data_1_0     (back_data_1_0),
    .in_valid_1_0    (back_valid_1_0),
    .in_ready_1_0    (back_ready_1_0),
    .in_data_1_1     (back_data_1_1),
    .in_valid_1_1    (back_valid_1_1),
    .in_ready_1_1    (back_ready_1_1),
    .in_data_1_2     (back_data_1_2),
    .in_valid_1_2    (back_valid_1_2),
    .in_ready_1_2    (back_ready_1_2),
    .in_data_1_3     (back_data_1_3),
    .in_valid_1_3    (back_valid_1_3),
    .in_ready_1_3    (back_ready_1_3),
    .in_data_1_4     (back_data_1_4),
    .in_valid_1_4    (back_valid_1_4),
    .in_ready_1_4    (back_ready_1_4),
    .in_data_1_5     (back_data_1_5),
    .in_valid_1_5    (back_valid_1_5),
    .in_ready_1_5    (back_ready_1_5),
    .in_data_1_6     (back_data_1_6),
    .in_valid_1_6    (back_valid_1_6),
    .in_ready_1_6    (back_ready_1_6),
    .in_data_1_7     (back_data_1_7),
    .in_valid_1_7    (back_valid_1_7),
    .in_ready_1_7    (back_ready_1_7),
    .in_data_1_8     (back_data_1_8),
    .in_valid_1_8    (back_valid_1_8),
    .in_ready_1_8    (back_ready_1_8),
    .in_data_1_9     (back_data_1_9),
    .in_valid_1_9    (back_valid_1_9),
    .in_ready_1_9    (back_ready_1_9),
    .in_data_1_10     (back_data_1_10),
    .in_valid_1_10    (back_valid_1_10),
    .in_ready_1_10    (back_ready_1_10),
    .in_data_1_11     (back_data_1_11),
    .in_valid_1_11    (back_valid_1_11),
    .in_ready_1_11    (back_ready_1_11),
    .in_data_1_12     (back_data_1_12),
    .in_valid_1_12    (back_valid_1_12),
    .in_ready_1_12    (back_ready_1_12),
    .in_data_1_13     (back_data_1_13),
    .in_valid_1_13    (back_valid_1_13),
    .in_ready_1_13    (back_ready_1_13),
    .in_data_1_14     (back_data_1_14),
    .in_valid_1_14    (back_valid_1_14),
    .in_ready_1_14    (back_ready_1_14),
    .in_data_1_15     (back_data_1_15),
    .in_valid_1_15    (back_valid_1_15),
    .in_ready_1_15    (back_ready_1_15),
    .in_data_1_16     (back_data_1_16),
    .in_valid_1_16    (back_valid_1_16),
    .in_ready_1_16    (back_ready_1_16),
    .in_data_1_17     (back_data_1_17),
    .in_valid_1_17    (back_valid_1_17),
    .in_ready_1_17    (back_ready_1_17),
    .in_data_1_18     (back_data_1_18),
    .in_valid_1_18    (back_valid_1_18),
    .in_ready_1_18    (back_ready_1_18),
    .in_data_1_19     (back_data_1_19),
    .in_valid_1_19    (back_valid_1_19),
    .in_ready_1_19    (back_ready_1_19),
    .in_data_1_20     (back_data_1_20),
    .in_valid_1_20    (back_valid_1_20),
    .in_ready_1_20    (back_ready_1_20),
    .in_data_1_21     (back_data_1_21),
    .in_valid_1_21    (back_valid_1_21),
    .in_ready_1_21    (back_ready_1_21),
    .in_data_1_22     (back_data_1_22),
    .in_valid_1_22    (back_valid_1_22),
    .in_ready_1_22    (back_ready_1_22),
    .in_data_1_23     (back_data_1_23),
    .in_valid_1_23    (back_valid_1_23),
    .in_ready_1_23    (back_ready_1_23),
    .in_data_1_24     (back_data_1_24),
    .in_valid_1_24    (back_valid_1_24),
    .in_ready_1_24    (back_ready_1_24),
    .in_data_1_25     (back_data_1_25),
    .in_valid_1_25    (back_valid_1_25),
    .in_ready_1_25    (back_ready_1_25),
    .in_data_1_26     (back_data_1_26),
    .in_valid_1_26    (back_valid_1_26),
    .in_ready_1_26    (back_ready_1_26),
    .in_data_1_27     (back_data_1_27),
    .in_valid_1_27    (back_valid_1_27),
    .in_ready_1_27    (back_ready_1_27),
    .in_data_1_28     (back_data_1_28),
    .in_valid_1_28    (back_valid_1_28),
    .in_ready_1_28    (back_ready_1_28),
    .in_data_1_29     (back_data_1_29),
    .in_valid_1_29    (back_valid_1_29),
    .in_ready_1_29    (back_ready_1_29),
    .in_data_1_30     (back_data_1_30),
    .in_valid_1_30    (back_valid_1_30),
    .in_ready_1_30    (back_ready_1_30),
    .in_data_1_31     (back_data_1_31),
    .in_valid_1_31    (back_valid_1_31),
    .in_ready_1_31    (back_ready_1_31),
    .in_data_2_0     (back_data_2_0),
    .in_valid_2_0    (back_valid_2_0),
    .in_ready_2_0    (back_ready_2_0),
    .in_data_2_1     (back_data_2_1),
    .in_valid_2_1    (back_valid_2_1),
    .in_ready_2_1    (back_ready_2_1),
    .in_data_2_2     (back_data_2_2),
    .in_valid_2_2    (back_valid_2_2),
    .in_ready_2_2    (back_ready_2_2),
    .in_data_2_3     (back_data_2_3),
    .in_valid_2_3    (back_valid_2_3),
    .in_ready_2_3    (back_ready_2_3),
    .in_data_2_4     (back_data_2_4),
    .in_valid_2_4    (back_valid_2_4),
    .in_ready_2_4    (back_ready_2_4),
    .in_data_2_5     (back_data_2_5),
    .in_valid_2_5    (back_valid_2_5),
    .in_ready_2_5    (back_ready_2_5),
    .in_data_2_6     (back_data_2_6),
    .in_valid_2_6    (back_valid_2_6),
    .in_ready_2_6    (back_ready_2_6),
    .in_data_2_7     (back_data_2_7),
    .in_valid_2_7    (back_valid_2_7),
    .in_ready_2_7    (back_ready_2_7),
    .in_data_2_8     (back_data_2_8),
    .in_valid_2_8    (back_valid_2_8),
    .in_ready_2_8    (back_ready_2_8),
    .in_data_2_9     (back_data_2_9),
    .in_valid_2_9    (back_valid_2_9),
    .in_ready_2_9    (back_ready_2_9),
    .in_data_2_10     (back_data_2_10),
    .in_valid_2_10    (back_valid_2_10),
    .in_ready_2_10    (back_ready_2_10),
    .in_data_2_11     (back_data_2_11),
    .in_valid_2_11    (back_valid_2_11),
    .in_ready_2_11    (back_ready_2_11),
    .in_data_2_12     (back_data_2_12),
    .in_valid_2_12    (back_valid_2_12),
    .in_ready_2_12    (back_ready_2_12),
    .in_data_2_13     (back_data_2_13),
    .in_valid_2_13    (back_valid_2_13),
    .in_ready_2_13    (back_ready_2_13),
    .in_data_2_14     (back_data_2_14),
    .in_valid_2_14    (back_valid_2_14),
    .in_ready_2_14    (back_ready_2_14),
    .in_data_2_15     (back_data_2_15),
    .in_valid_2_15    (back_valid_2_15),
    .in_ready_2_15    (back_ready_2_15),
    .in_data_2_16     (back_data_2_16),
    .in_valid_2_16    (back_valid_2_16),
    .in_ready_2_16    (back_ready_2_16),
    .in_data_2_17     (back_data_2_17),
    .in_valid_2_17    (back_valid_2_17),
    .in_ready_2_17    (back_ready_2_17),
    .in_data_2_18     (back_data_2_18),
    .in_valid_2_18    (back_valid_2_18),
    .in_ready_2_18    (back_ready_2_18),
    .in_data_2_19     (back_data_2_19),
    .in_valid_2_19    (back_valid_2_19),
    .in_ready_2_19    (back_ready_2_19),
    .in_data_2_20     (back_data_2_20),
    .in_valid_2_20    (back_valid_2_20),
    .in_ready_2_20    (back_ready_2_20),
    .in_data_2_21     (back_data_2_21),
    .in_valid_2_21    (back_valid_2_21),
    .in_ready_2_21    (back_ready_2_21),
    .in_data_2_22     (back_data_2_22),
    .in_valid_2_22    (back_valid_2_22),
    .in_ready_2_22    (back_ready_2_22),
    .in_data_2_23     (back_data_2_23),
    .in_valid_2_23    (back_valid_2_23),
    .in_ready_2_23    (back_ready_2_23),
    .in_data_2_24     (back_data_2_24),
    .in_valid_2_24    (back_valid_2_24),
    .in_ready_2_24    (back_ready_2_24),
    .in_data_2_25     (back_data_2_25),
    .in_valid_2_25    (back_valid_2_25),
    .in_ready_2_25    (back_ready_2_25),
    .in_data_2_26     (back_data_2_26),
    .in_valid_2_26    (back_valid_2_26),
    .in_ready_2_26    (back_ready_2_26),
    .in_data_2_27     (back_data_2_27),
    .in_valid_2_27    (back_valid_2_27),
    .in_ready_2_27    (back_ready_2_27),
    .in_data_2_28     (back_data_2_28),
    .in_valid_2_28    (back_valid_2_28),
    .in_ready_2_28    (back_ready_2_28),
    .in_data_2_29     (back_data_2_29),
    .in_valid_2_29    (back_valid_2_29),
    .in_ready_2_29    (back_ready_2_29),
    .in_data_2_30     (back_data_2_30),
    .in_valid_2_30    (back_valid_2_30),
    .in_ready_2_30    (back_ready_2_30),
    .in_data_2_31     (back_data_2_31),
    .in_valid_2_31    (back_valid_2_31),
    .in_ready_2_31    (back_ready_2_31),
    .in_data_3_0     (back_data_3_0),
    .in_valid_3_0    (back_valid_3_0),
    .in_ready_3_0    (back_ready_3_0),
    .in_data_3_1     (back_data_3_1),
    .in_valid_3_1    (back_valid_3_1),
    .in_ready_3_1    (back_ready_3_1),
    .in_data_3_2     (back_data_3_2),
    .in_valid_3_2    (back_valid_3_2),
    .in_ready_3_2    (back_ready_3_2),
    .in_data_3_3     (back_data_3_3),
    .in_valid_3_3    (back_valid_3_3),
    .in_ready_3_3    (back_ready_3_3),
    .in_data_3_4     (back_data_3_4),
    .in_valid_3_4    (back_valid_3_4),
    .in_ready_3_4    (back_ready_3_4),
    .in_data_3_5     (back_data_3_5),
    .in_valid_3_5    (back_valid_3_5),
    .in_ready_3_5    (back_ready_3_5),
    .in_data_3_6     (back_data_3_6),
    .in_valid_3_6    (back_valid_3_6),
    .in_ready_3_6    (back_ready_3_6),
    .in_data_3_7     (back_data_3_7),
    .in_valid_3_7    (back_valid_3_7),
    .in_ready_3_7    (back_ready_3_7),
    .in_data_3_8     (back_data_3_8),
    .in_valid_3_8    (back_valid_3_8),
    .in_ready_3_8    (back_ready_3_8),
    .in_data_3_9     (back_data_3_9),
    .in_valid_3_9    (back_valid_3_9),
    .in_ready_3_9    (back_ready_3_9),
    .in_data_3_10     (back_data_3_10),
    .in_valid_3_10    (back_valid_3_10),
    .in_ready_3_10    (back_ready_3_10),
    .in_data_3_11     (back_data_3_11),
    .in_valid_3_11    (back_valid_3_11),
    .in_ready_3_11    (back_ready_3_11),
    .in_data_3_12     (back_data_3_12),
    .in_valid_3_12    (back_valid_3_12),
    .in_ready_3_12    (back_ready_3_12),
    .in_data_3_13     (back_data_3_13),
    .in_valid_3_13    (back_valid_3_13),
    .in_ready_3_13    (back_ready_3_13),
    .in_data_3_14     (back_data_3_14),
    .in_valid_3_14    (back_valid_3_14),
    .in_ready_3_14    (back_ready_3_14),
    .in_data_3_15     (back_data_3_15),
    .in_valid_3_15    (back_valid_3_15),
    .in_ready_3_15    (back_ready_3_15),
    .in_data_3_16     (back_data_3_16),
    .in_valid_3_16    (back_valid_3_16),
    .in_ready_3_16    (back_ready_3_16),
    .in_data_3_17     (back_data_3_17),
    .in_valid_3_17    (back_valid_3_17),
    .in_ready_3_17    (back_ready_3_17),
    .in_data_3_18     (back_data_3_18),
    .in_valid_3_18    (back_valid_3_18),
    .in_ready_3_18    (back_ready_3_18),
    .in_data_3_19     (back_data_3_19),
    .in_valid_3_19    (back_valid_3_19),
    .in_ready_3_19    (back_ready_3_19),
    .in_data_3_20     (back_data_3_20),
    .in_valid_3_20    (back_valid_3_20),
    .in_ready_3_20    (back_ready_3_20),
    .in_data_3_21     (back_data_3_21),
    .in_valid_3_21    (back_valid_3_21),
    .in_ready_3_21    (back_ready_3_21),
    .in_data_3_22     (back_data_3_22),
    .in_valid_3_22    (back_valid_3_22),
    .in_ready_3_22    (back_ready_3_22),
    .in_data_3_23     (back_data_3_23),
    .in_valid_3_23    (back_valid_3_23),
    .in_ready_3_23    (back_ready_3_23),
    .in_data_3_24     (back_data_3_24),
    .in_valid_3_24    (back_valid_3_24),
    .in_ready_3_24    (back_ready_3_24),
    .in_data_3_25     (back_data_3_25),
    .in_valid_3_25    (back_valid_3_25),
    .in_ready_3_25    (back_ready_3_25),
    .in_data_3_26     (back_data_3_26),
    .in_valid_3_26    (back_valid_3_26),
    .in_ready_3_26    (back_ready_3_26),
    .in_data_3_27     (back_data_3_27),
    .in_valid_3_27    (back_valid_3_27),
    .in_ready_3_27    (back_ready_3_27),
    .in_data_3_28     (back_data_3_28),
    .in_valid_3_28    (back_valid_3_28),
    .in_ready_3_28    (back_ready_3_28),
    .in_data_3_29     (back_data_3_29),
    .in_valid_3_29    (back_valid_3_29),
    .in_ready_3_29    (back_ready_3_29),
    .in_data_3_30     (back_data_3_30),
    .in_valid_3_30    (back_valid_3_30),
    .in_ready_3_30    (back_ready_3_30),
    .in_data_3_31     (back_data_3_31),
    .in_valid_3_31    (back_valid_3_31),
    .in_ready_3_31    (back_ready_3_31),
    .in_data_4_0     (back_data_4_0),
    .in_valid_4_0    (back_valid_4_0),
    .in_ready_4_0    (back_ready_4_0),
    .in_data_4_1     (back_data_4_1),
    .in_valid_4_1    (back_valid_4_1),
    .in_ready_4_1    (back_ready_4_1),
    .in_data_4_2     (back_data_4_2),
    .in_valid_4_2    (back_valid_4_2),
    .in_ready_4_2    (back_ready_4_2),
    .in_data_4_3     (back_data_4_3),
    .in_valid_4_3    (back_valid_4_3),
    .in_ready_4_3    (back_ready_4_3),
    .in_data_4_4     (back_data_4_4),
    .in_valid_4_4    (back_valid_4_4),
    .in_ready_4_4    (back_ready_4_4),
    .in_data_4_5     (back_data_4_5),
    .in_valid_4_5    (back_valid_4_5),
    .in_ready_4_5    (back_ready_4_5),
    .in_data_4_6     (back_data_4_6),
    .in_valid_4_6    (back_valid_4_6),
    .in_ready_4_6    (back_ready_4_6),
    .in_data_4_7     (back_data_4_7),
    .in_valid_4_7    (back_valid_4_7),
    .in_ready_4_7    (back_ready_4_7),
    .in_data_4_8     (back_data_4_8),
    .in_valid_4_8    (back_valid_4_8),
    .in_ready_4_8    (back_ready_4_8),
    .in_data_4_9     (back_data_4_9),
    .in_valid_4_9    (back_valid_4_9),
    .in_ready_4_9    (back_ready_4_9),
    .in_data_4_10     (back_data_4_10),
    .in_valid_4_10    (back_valid_4_10),
    .in_ready_4_10    (back_ready_4_10),
    .in_data_4_11     (back_data_4_11),
    .in_valid_4_11    (back_valid_4_11),
    .in_ready_4_11    (back_ready_4_11),
    .in_data_4_12     (back_data_4_12),
    .in_valid_4_12    (back_valid_4_12),
    .in_ready_4_12    (back_ready_4_12),
    .in_data_4_13     (back_data_4_13),
    .in_valid_4_13    (back_valid_4_13),
    .in_ready_4_13    (back_ready_4_13),
    .in_data_4_14     (back_data_4_14),
    .in_valid_4_14    (back_valid_4_14),
    .in_ready_4_14    (back_ready_4_14),
    .in_data_4_15     (back_data_4_15),
    .in_valid_4_15    (back_valid_4_15),
    .in_ready_4_15    (back_ready_4_15),
    .in_data_4_16     (back_data_4_16),
    .in_valid_4_16    (back_valid_4_16),
    .in_ready_4_16    (back_ready_4_16),
    .in_data_4_17     (back_data_4_17),
    .in_valid_4_17    (back_valid_4_17),
    .in_ready_4_17    (back_ready_4_17),
    .in_data_4_18     (back_data_4_18),
    .in_valid_4_18    (back_valid_4_18),
    .in_ready_4_18    (back_ready_4_18),
    .in_data_4_19     (back_data_4_19),
    .in_valid_4_19    (back_valid_4_19),
    .in_ready_4_19    (back_ready_4_19),
    .in_data_4_20     (back_data_4_20),
    .in_valid_4_20    (back_valid_4_20),
    .in_ready_4_20    (back_ready_4_20),
    .in_data_4_21     (back_data_4_21),
    .in_valid_4_21    (back_valid_4_21),
    .in_ready_4_21    (back_ready_4_21),
    .in_data_4_22     (back_data_4_22),
    .in_valid_4_22    (back_valid_4_22),
    .in_ready_4_22    (back_ready_4_22),
    .in_data_4_23     (back_data_4_23),
    .in_valid_4_23    (back_valid_4_23),
    .in_ready_4_23    (back_ready_4_23),
    .in_data_4_24     (back_data_4_24),
    .in_valid_4_24    (back_valid_4_24),
    .in_ready_4_24    (back_ready_4_24),
    .in_data_4_25     (back_data_4_25),
    .in_valid_4_25    (back_valid_4_25),
    .in_ready_4_25    (back_ready_4_25),
    .in_data_4_26     (back_data_4_26),
    .in_valid_4_26    (back_valid_4_26),
    .in_ready_4_26    (back_ready_4_26),
    .in_data_4_27     (back_data_4_27),
    .in_valid_4_27    (back_valid_4_27),
    .in_ready_4_27    (back_ready_4_27),
    .in_data_4_28     (back_data_4_28),
    .in_valid_4_28    (back_valid_4_28),
    .in_ready_4_28    (back_ready_4_28),
    .in_data_4_29     (back_data_4_29),
    .in_valid_4_29    (back_valid_4_29),
    .in_ready_4_29    (back_ready_4_29),
    .in_data_4_30     (back_data_4_30),
    .in_valid_4_30    (back_valid_4_30),
    .in_ready_4_30    (back_ready_4_30),
    .in_data_4_31     (back_data_4_31),
    .in_valid_4_31    (back_valid_4_31),
    .in_ready_4_31    (back_ready_4_31),
    .in_data_5_0     (back_data_5_0),
    .in_valid_5_0    (back_valid_5_0),
    .in_ready_5_0    (back_ready_5_0),
    .in_data_5_1     (back_data_5_1),
    .in_valid_5_1    (back_valid_5_1),
    .in_ready_5_1    (back_ready_5_1),
    .in_data_5_2     (back_data_5_2),
    .in_valid_5_2    (back_valid_5_2),
    .in_ready_5_2    (back_ready_5_2),
    .in_data_5_3     (back_data_5_3),
    .in_valid_5_3    (back_valid_5_3),
    .in_ready_5_3    (back_ready_5_3),
    .in_data_5_4     (back_data_5_4),
    .in_valid_5_4    (back_valid_5_4),
    .in_ready_5_4    (back_ready_5_4),
    .in_data_5_5     (back_data_5_5),
    .in_valid_5_5    (back_valid_5_5),
    .in_ready_5_5    (back_ready_5_5),
    .in_data_5_6     (back_data_5_6),
    .in_valid_5_6    (back_valid_5_6),
    .in_ready_5_6    (back_ready_5_6),
    .in_data_5_7     (back_data_5_7),
    .in_valid_5_7    (back_valid_5_7),
    .in_ready_5_7    (back_ready_5_7),
    .in_data_5_8     (back_data_5_8),
    .in_valid_5_8    (back_valid_5_8),
    .in_ready_5_8    (back_ready_5_8),
    .in_data_5_9     (back_data_5_9),
    .in_valid_5_9    (back_valid_5_9),
    .in_ready_5_9    (back_ready_5_9),
    .in_data_5_10     (back_data_5_10),
    .in_valid_5_10    (back_valid_5_10),
    .in_ready_5_10    (back_ready_5_10),
    .in_data_5_11     (back_data_5_11),
    .in_valid_5_11    (back_valid_5_11),
    .in_ready_5_11    (back_ready_5_11),
    .in_data_5_12     (back_data_5_12),
    .in_valid_5_12    (back_valid_5_12),
    .in_ready_5_12    (back_ready_5_12),
    .in_data_5_13     (back_data_5_13),
    .in_valid_5_13    (back_valid_5_13),
    .in_ready_5_13    (back_ready_5_13),
    .in_data_5_14     (back_data_5_14),
    .in_valid_5_14    (back_valid_5_14),
    .in_ready_5_14    (back_ready_5_14),
    .in_data_5_15     (back_data_5_15),
    .in_valid_5_15    (back_valid_5_15),
    .in_ready_5_15    (back_ready_5_15),
    .in_data_5_16     (back_data_5_16),
    .in_valid_5_16    (back_valid_5_16),
    .in_ready_5_16    (back_ready_5_16),
    .in_data_5_17     (back_data_5_17),
    .in_valid_5_17    (back_valid_5_17),
    .in_ready_5_17    (back_ready_5_17),
    .in_data_5_18     (back_data_5_18),
    .in_valid_5_18    (back_valid_5_18),
    .in_ready_5_18    (back_ready_5_18),
    .in_data_5_19     (back_data_5_19),
    .in_valid_5_19    (back_valid_5_19),
    .in_ready_5_19    (back_ready_5_19),
    .in_data_5_20     (back_data_5_20),
    .in_valid_5_20    (back_valid_5_20),
    .in_ready_5_20    (back_ready_5_20),
    .in_data_5_21     (back_data_5_21),
    .in_valid_5_21    (back_valid_5_21),
    .in_ready_5_21    (back_ready_5_21),
    .in_data_5_22     (back_data_5_22),
    .in_valid_5_22    (back_valid_5_22),
    .in_ready_5_22    (back_ready_5_22),
    .in_data_5_23     (back_data_5_23),
    .in_valid_5_23    (back_valid_5_23),
    .in_ready_5_23    (back_ready_5_23),
    .in_data_5_24     (back_data_5_24),
    .in_valid_5_24    (back_valid_5_24),
    .in_ready_5_24    (back_ready_5_24),
    .in_data_5_25     (back_data_5_25),
    .in_valid_5_25    (back_valid_5_25),
    .in_ready_5_25    (back_ready_5_25),
    .in_data_5_26     (back_data_5_26),
    .in_valid_5_26    (back_valid_5_26),
    .in_ready_5_26    (back_ready_5_26),
    .in_data_5_27     (back_data_5_27),
    .in_valid_5_27    (back_valid_5_27),
    .in_ready_5_27    (back_ready_5_27),
    .in_data_5_28     (back_data_5_28),
    .in_valid_5_28    (back_valid_5_28),
    .in_ready_5_28    (back_ready_5_28),
    .in_data_5_29     (back_data_5_29),
    .in_valid_5_29    (back_valid_5_29),
    .in_ready_5_29    (back_ready_5_29),
    .in_data_5_30     (back_data_5_30),
    .in_valid_5_30    (back_valid_5_30),
    .in_ready_5_30    (back_ready_5_30),
    .in_data_5_31     (back_data_5_31),
    .in_valid_5_31    (back_valid_5_31),
    .in_ready_5_31    (back_ready_5_31),
    .in_data_6_0     (back_data_6_0),
    .in_valid_6_0    (back_valid_6_0),
    .in_ready_6_0    (back_ready_6_0),
    .in_data_6_1     (back_data_6_1),
    .in_valid_6_1    (back_valid_6_1),
    .in_ready_6_1    (back_ready_6_1),
    .in_data_6_2     (back_data_6_2),
    .in_valid_6_2    (back_valid_6_2),
    .in_ready_6_2    (back_ready_6_2),
    .in_data_6_3     (back_data_6_3),
    .in_valid_6_3    (back_valid_6_3),
    .in_ready_6_3    (back_ready_6_3),
    .in_data_6_4     (back_data_6_4),
    .in_valid_6_4    (back_valid_6_4),
    .in_ready_6_4    (back_ready_6_4),
    .in_data_6_5     (back_data_6_5),
    .in_valid_6_5    (back_valid_6_5),
    .in_ready_6_5    (back_ready_6_5),
    .in_data_6_6     (back_data_6_6),
    .in_valid_6_6    (back_valid_6_6),
    .in_ready_6_6    (back_ready_6_6),
    .in_data_6_7     (back_data_6_7),
    .in_valid_6_7    (back_valid_6_7),
    .in_ready_6_7    (back_ready_6_7),
    .in_data_6_8     (back_data_6_8),
    .in_valid_6_8    (back_valid_6_8),
    .in_ready_6_8    (back_ready_6_8),
    .in_data_6_9     (back_data_6_9),
    .in_valid_6_9    (back_valid_6_9),
    .in_ready_6_9    (back_ready_6_9),
    .in_data_6_10     (back_data_6_10),
    .in_valid_6_10    (back_valid_6_10),
    .in_ready_6_10    (back_ready_6_10),
    .in_data_6_11     (back_data_6_11),
    .in_valid_6_11    (back_valid_6_11),
    .in_ready_6_11    (back_ready_6_11),
    .in_data_6_12     (back_data_6_12),
    .in_valid_6_12    (back_valid_6_12),
    .in_ready_6_12    (back_ready_6_12),
    .in_data_6_13     (back_data_6_13),
    .in_valid_6_13    (back_valid_6_13),
    .in_ready_6_13    (back_ready_6_13),
    .in_data_6_14     (back_data_6_14),
    .in_valid_6_14    (back_valid_6_14),
    .in_ready_6_14    (back_ready_6_14),
    .in_data_6_15     (back_data_6_15),
    .in_valid_6_15    (back_valid_6_15),
    .in_ready_6_15    (back_ready_6_15),
    .in_data_6_16     (back_data_6_16),
    .in_valid_6_16    (back_valid_6_16),
    .in_ready_6_16    (back_ready_6_16),
    .in_data_6_17     (back_data_6_17),
    .in_valid_6_17    (back_valid_6_17),
    .in_ready_6_17    (back_ready_6_17),
    .in_data_6_18     (back_data_6_18),
    .in_valid_6_18    (back_valid_6_18),
    .in_ready_6_18    (back_ready_6_18),
    .in_data_6_19     (back_data_6_19),
    .in_valid_6_19    (back_valid_6_19),
    .in_ready_6_19    (back_ready_6_19),
    .in_data_6_20     (back_data_6_20),
    .in_valid_6_20    (back_valid_6_20),
    .in_ready_6_20    (back_ready_6_20),
    .in_data_6_21     (back_data_6_21),
    .in_valid_6_21    (back_valid_6_21),
    .in_ready_6_21    (back_ready_6_21),
    .in_data_6_22     (back_data_6_22),
    .in_valid_6_22    (back_valid_6_22),
    .in_ready_6_22    (back_ready_6_22),
    .in_data_6_23     (back_data_6_23),
    .in_valid_6_23    (back_valid_6_23),
    .in_ready_6_23    (back_ready_6_23),
    .in_data_6_24     (back_data_6_24),
    .in_valid_6_24    (back_valid_6_24),
    .in_ready_6_24    (back_ready_6_24),
    .in_data_6_25     (back_data_6_25),
    .in_valid_6_25    (back_valid_6_25),
    .in_ready_6_25    (back_ready_6_25),
    .in_data_6_26     (back_data_6_26),
    .in_valid_6_26    (back_valid_6_26),
    .in_ready_6_26    (back_ready_6_26),
    .in_data_6_27     (back_data_6_27),
    .in_valid_6_27    (back_valid_6_27),
    .in_ready_6_27    (back_ready_6_27),
    .in_data_6_28     (back_data_6_28),
    .in_valid_6_28    (back_valid_6_28),
    .in_ready_6_28    (back_ready_6_28),
    .in_data_6_29     (back_data_6_29),
    .in_valid_6_29    (back_valid_6_29),
    .in_ready_6_29    (back_ready_6_29),
    .in_data_6_30     (back_data_6_30),
    .in_valid_6_30    (back_valid_6_30),
    .in_ready_6_30    (back_ready_6_30),
    .in_data_6_31     (back_data_6_31),
    .in_valid_6_31    (back_valid_6_31),
    .in_ready_6_31    (back_ready_6_31),
    .in_data_7_0     (back_data_7_0),
    .in_valid_7_0    (back_valid_7_0),
    .in_ready_7_0    (back_ready_7_0),
    .in_data_7_1     (back_data_7_1),
    .in_valid_7_1    (back_valid_7_1),
    .in_ready_7_1    (back_ready_7_1),
    .in_data_7_2     (back_data_7_2),
    .in_valid_7_2    (back_valid_7_2),
    .in_ready_7_2    (back_ready_7_2),
    .in_data_7_3     (back_data_7_3),
    .in_valid_7_3    (back_valid_7_3),
    .in_ready_7_3    (back_ready_7_3),
    .in_data_7_4     (back_data_7_4),
    .in_valid_7_4    (back_valid_7_4),
    .in_ready_7_4    (back_ready_7_4),
    .in_data_7_5     (back_data_7_5),
    .in_valid_7_5    (back_valid_7_5),
    .in_ready_7_5    (back_ready_7_5),
    .in_data_7_6     (back_data_7_6),
    .in_valid_7_6    (back_valid_7_6),
    .in_ready_7_6    (back_ready_7_6),
    .in_data_7_7     (back_data_7_7),
    .in_valid_7_7    (back_valid_7_7),
    .in_ready_7_7    (back_ready_7_7),
    .in_data_7_8     (back_data_7_8),
    .in_valid_7_8    (back_valid_7_8),
    .in_ready_7_8    (back_ready_7_8),
    .in_data_7_9     (back_data_7_9),
    .in_valid_7_9    (back_valid_7_9),
    .in_ready_7_9    (back_ready_7_9),
    .in_data_7_10     (back_data_7_10),
    .in_valid_7_10    (back_valid_7_10),
    .in_ready_7_10    (back_ready_7_10),
    .in_data_7_11     (back_data_7_11),
    .in_valid_7_11    (back_valid_7_11),
    .in_ready_7_11    (back_ready_7_11),
    .in_data_7_12     (back_data_7_12),
    .in_valid_7_12    (back_valid_7_12),
    .in_ready_7_12    (back_ready_7_12),
    .in_data_7_13     (back_data_7_13),
    .in_valid_7_13    (back_valid_7_13),
    .in_ready_7_13    (back_ready_7_13),
    .in_data_7_14     (back_data_7_14),
    .in_valid_7_14    (back_valid_7_14),
    .in_ready_7_14    (back_ready_7_14),
    .in_data_7_15     (back_data_7_15),
    .in_valid_7_15    (back_valid_7_15),
    .in_ready_7_15    (back_ready_7_15),
    .in_data_7_16     (back_data_7_16),
    .in_valid_7_16    (back_valid_7_16),
    .in_ready_7_16    (back_ready_7_16),
    .in_data_7_17     (back_data_7_17),
    .in_valid_7_17    (back_valid_7_17),
    .in_ready_7_17    (back_ready_7_17),
    .in_data_7_18     (back_data_7_18),
    .in_valid_7_18    (back_valid_7_18),
    .in_ready_7_18    (back_ready_7_18),
    .in_data_7_19     (back_data_7_19),
    .in_valid_7_19    (back_valid_7_19),
    .in_ready_7_19    (back_ready_7_19),
    .in_data_7_20     (back_data_7_20),
    .in_valid_7_20    (back_valid_7_20),
    .in_ready_7_20    (back_ready_7_20),
    .in_data_7_21     (back_data_7_21),
    .in_valid_7_21    (back_valid_7_21),
    .in_ready_7_21    (back_ready_7_21),
    .in_data_7_22     (back_data_7_22),
    .in_valid_7_22    (back_valid_7_22),
    .in_ready_7_22    (back_ready_7_22),
    .in_data_7_23     (back_data_7_23),
    .in_valid_7_23    (back_valid_7_23),
    .in_ready_7_23    (back_ready_7_23),
    .in_data_7_24     (back_data_7_24),
    .in_valid_7_24    (back_valid_7_24),
    .in_ready_7_24    (back_ready_7_24),
    .in_data_7_25     (back_data_7_25),
    .in_valid_7_25    (back_valid_7_25),
    .in_ready_7_25    (back_ready_7_25),
    .in_data_7_26     (back_data_7_26),
    .in_valid_7_26    (back_valid_7_26),
    .in_ready_7_26    (back_ready_7_26),
    .in_data_7_27     (back_data_7_27),
    .in_valid_7_27    (back_valid_7_27),
    .in_ready_7_27    (back_ready_7_27),
    .in_data_7_28     (back_data_7_28),
    .in_valid_7_28    (back_valid_7_28),
    .in_ready_7_28    (back_ready_7_28),
    .in_data_7_29     (back_data_7_29),
    .in_valid_7_29    (back_valid_7_29),
    .in_ready_7_29    (back_ready_7_29),
    .in_data_7_30     (back_data_7_30),
    .in_valid_7_30    (back_valid_7_30),
    .in_ready_7_30    (back_ready_7_30),
    .in_data_7_31     (back_data_7_31),
    .in_valid_7_31    (back_valid_7_31),
    .in_ready_7_31    (back_ready_7_31),
    .out_usr_data            (out_usr_data),
    .out_usr_valid           (out_usr_valid),
    .out_usr_sop             (out_usr_sop),
    .out_usr_eop             (out_usr_eop),
    .out_usr_empty           (out_usr_empty),
    .out_usr_ready           (out_usr_ready)
);


//Cross clock domain
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_0"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_0 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_0_r2),              
    .in_valid          (din_valid_0_0_r2),             
    .in_ready          (din_ready_0_0),             
    .out_data          (back_data_0_0),              
    .out_valid         (back_valid_0_0),             
    .out_ready         (back_ready_0_0),             
    .fill_level        (din_csr_readdata_0_0),
    .almost_full       (din_almost_full_0_0),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_1"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_1 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_1_r2),              
    .in_valid          (din_valid_0_1_r2),             
    .in_ready          (din_ready_0_1),             
    .out_data          (back_data_0_1),              
    .out_valid         (back_valid_0_1),             
    .out_ready         (back_ready_0_1),             
    .fill_level        (din_csr_readdata_0_1),
    .almost_full       (din_almost_full_0_1),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_2"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_2 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_2_r2),              
    .in_valid          (din_valid_0_2_r2),             
    .in_ready          (din_ready_0_2),             
    .out_data          (back_data_0_2),              
    .out_valid         (back_valid_0_2),             
    .out_ready         (back_ready_0_2),             
    .fill_level        (din_csr_readdata_0_2),
    .almost_full       (din_almost_full_0_2),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_3"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_3 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_3_r2),              
    .in_valid          (din_valid_0_3_r2),             
    .in_ready          (din_ready_0_3),             
    .out_data          (back_data_0_3),              
    .out_valid         (back_valid_0_3),             
    .out_ready         (back_ready_0_3),             
    .fill_level        (din_csr_readdata_0_3),
    .almost_full       (din_almost_full_0_3),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_4"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_4 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_4_r2),              
    .in_valid          (din_valid_0_4_r2),             
    .in_ready          (din_ready_0_4),             
    .out_data          (back_data_0_4),              
    .out_valid         (back_valid_0_4),             
    .out_ready         (back_ready_0_4),             
    .fill_level        (din_csr_readdata_0_4),
    .almost_full       (din_almost_full_0_4),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_5"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_5 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_5_r2),              
    .in_valid          (din_valid_0_5_r2),             
    .in_ready          (din_ready_0_5),             
    .out_data          (back_data_0_5),              
    .out_valid         (back_valid_0_5),             
    .out_ready         (back_ready_0_5),             
    .fill_level        (din_csr_readdata_0_5),
    .almost_full       (din_almost_full_0_5),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_6"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_6 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_6_r2),              
    .in_valid          (din_valid_0_6_r2),             
    .in_ready          (din_ready_0_6),             
    .out_data          (back_data_0_6),              
    .out_valid         (back_valid_0_6),             
    .out_ready         (back_ready_0_6),             
    .fill_level        (din_csr_readdata_0_6),
    .almost_full       (din_almost_full_0_6),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_7"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_7 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_7_r2),              
    .in_valid          (din_valid_0_7_r2),             
    .in_ready          (din_ready_0_7),             
    .out_data          (back_data_0_7),              
    .out_valid         (back_valid_0_7),             
    .out_ready         (back_ready_0_7),             
    .fill_level        (din_csr_readdata_0_7),
    .almost_full       (din_almost_full_0_7),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_8"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_8 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_8_r2),              
    .in_valid          (din_valid_0_8_r2),             
    .in_ready          (din_ready_0_8),             
    .out_data          (back_data_0_8),              
    .out_valid         (back_valid_0_8),             
    .out_ready         (back_ready_0_8),             
    .fill_level        (din_csr_readdata_0_8),
    .almost_full       (din_almost_full_0_8),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_9"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_9 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_9_r2),              
    .in_valid          (din_valid_0_9_r2),             
    .in_ready          (din_ready_0_9),             
    .out_data          (back_data_0_9),              
    .out_valid         (back_valid_0_9),             
    .out_ready         (back_ready_0_9),             
    .fill_level        (din_csr_readdata_0_9),
    .almost_full       (din_almost_full_0_9),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_10"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_10 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_10_r2),              
    .in_valid          (din_valid_0_10_r2),             
    .in_ready          (din_ready_0_10),             
    .out_data          (back_data_0_10),              
    .out_valid         (back_valid_0_10),             
    .out_ready         (back_ready_0_10),             
    .fill_level        (din_csr_readdata_0_10),
    .almost_full       (din_almost_full_0_10),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_11"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_11 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_11_r2),              
    .in_valid          (din_valid_0_11_r2),             
    .in_ready          (din_ready_0_11),             
    .out_data          (back_data_0_11),              
    .out_valid         (back_valid_0_11),             
    .out_ready         (back_ready_0_11),             
    .fill_level        (din_csr_readdata_0_11),
    .almost_full       (din_almost_full_0_11),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_12"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_12 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_12_r2),              
    .in_valid          (din_valid_0_12_r2),             
    .in_ready          (din_ready_0_12),             
    .out_data          (back_data_0_12),              
    .out_valid         (back_valid_0_12),             
    .out_ready         (back_ready_0_12),             
    .fill_level        (din_csr_readdata_0_12),
    .almost_full       (din_almost_full_0_12),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_13"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_13 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_13_r2),              
    .in_valid          (din_valid_0_13_r2),             
    .in_ready          (din_ready_0_13),             
    .out_data          (back_data_0_13),              
    .out_valid         (back_valid_0_13),             
    .out_ready         (back_ready_0_13),             
    .fill_level        (din_csr_readdata_0_13),
    .almost_full       (din_almost_full_0_13),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_14"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_14 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_14_r2),              
    .in_valid          (din_valid_0_14_r2),             
    .in_ready          (din_ready_0_14),             
    .out_data          (back_data_0_14),              
    .out_valid         (back_valid_0_14),             
    .out_ready         (back_ready_0_14),             
    .fill_level        (din_csr_readdata_0_14),
    .almost_full       (din_almost_full_0_14),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_15"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_15 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_15_r2),              
    .in_valid          (din_valid_0_15_r2),             
    .in_ready          (din_ready_0_15),             
    .out_data          (back_data_0_15),              
    .out_valid         (back_valid_0_15),             
    .out_ready         (back_ready_0_15),             
    .fill_level        (din_csr_readdata_0_15),
    .almost_full       (din_almost_full_0_15),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_16"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_16 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_16_r2),              
    .in_valid          (din_valid_0_16_r2),             
    .in_ready          (din_ready_0_16),             
    .out_data          (back_data_0_16),              
    .out_valid         (back_valid_0_16),             
    .out_ready         (back_ready_0_16),             
    .fill_level        (din_csr_readdata_0_16),
    .almost_full       (din_almost_full_0_16),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_17"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_17 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_17_r2),              
    .in_valid          (din_valid_0_17_r2),             
    .in_ready          (din_ready_0_17),             
    .out_data          (back_data_0_17),              
    .out_valid         (back_valid_0_17),             
    .out_ready         (back_ready_0_17),             
    .fill_level        (din_csr_readdata_0_17),
    .almost_full       (din_almost_full_0_17),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_18"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_18 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_18_r2),              
    .in_valid          (din_valid_0_18_r2),             
    .in_ready          (din_ready_0_18),             
    .out_data          (back_data_0_18),              
    .out_valid         (back_valid_0_18),             
    .out_ready         (back_ready_0_18),             
    .fill_level        (din_csr_readdata_0_18),
    .almost_full       (din_almost_full_0_18),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_19"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_19 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_19_r2),              
    .in_valid          (din_valid_0_19_r2),             
    .in_ready          (din_ready_0_19),             
    .out_data          (back_data_0_19),              
    .out_valid         (back_valid_0_19),             
    .out_ready         (back_ready_0_19),             
    .fill_level        (din_csr_readdata_0_19),
    .almost_full       (din_almost_full_0_19),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_20"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_20 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_20_r2),              
    .in_valid          (din_valid_0_20_r2),             
    .in_ready          (din_ready_0_20),             
    .out_data          (back_data_0_20),              
    .out_valid         (back_valid_0_20),             
    .out_ready         (back_ready_0_20),             
    .fill_level        (din_csr_readdata_0_20),
    .almost_full       (din_almost_full_0_20),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_21"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_21 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_21_r2),              
    .in_valid          (din_valid_0_21_r2),             
    .in_ready          (din_ready_0_21),             
    .out_data          (back_data_0_21),              
    .out_valid         (back_valid_0_21),             
    .out_ready         (back_ready_0_21),             
    .fill_level        (din_csr_readdata_0_21),
    .almost_full       (din_almost_full_0_21),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_22"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_22 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_22_r2),              
    .in_valid          (din_valid_0_22_r2),             
    .in_ready          (din_ready_0_22),             
    .out_data          (back_data_0_22),              
    .out_valid         (back_valid_0_22),             
    .out_ready         (back_ready_0_22),             
    .fill_level        (din_csr_readdata_0_22),
    .almost_full       (din_almost_full_0_22),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_23"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_23 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_23_r2),              
    .in_valid          (din_valid_0_23_r2),             
    .in_ready          (din_ready_0_23),             
    .out_data          (back_data_0_23),              
    .out_valid         (back_valid_0_23),             
    .out_ready         (back_ready_0_23),             
    .fill_level        (din_csr_readdata_0_23),
    .almost_full       (din_almost_full_0_23),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_24"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_24 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_24_r2),              
    .in_valid          (din_valid_0_24_r2),             
    .in_ready          (din_ready_0_24),             
    .out_data          (back_data_0_24),              
    .out_valid         (back_valid_0_24),             
    .out_ready         (back_ready_0_24),             
    .fill_level        (din_csr_readdata_0_24),
    .almost_full       (din_almost_full_0_24),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_25"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_25 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_25_r2),              
    .in_valid          (din_valid_0_25_r2),             
    .in_ready          (din_ready_0_25),             
    .out_data          (back_data_0_25),              
    .out_valid         (back_valid_0_25),             
    .out_ready         (back_ready_0_25),             
    .fill_level        (din_csr_readdata_0_25),
    .almost_full       (din_almost_full_0_25),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_26"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_26 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_26_r2),              
    .in_valid          (din_valid_0_26_r2),             
    .in_ready          (din_ready_0_26),             
    .out_data          (back_data_0_26),              
    .out_valid         (back_valid_0_26),             
    .out_ready         (back_ready_0_26),             
    .fill_level        (din_csr_readdata_0_26),
    .almost_full       (din_almost_full_0_26),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_27"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_27 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_27_r2),              
    .in_valid          (din_valid_0_27_r2),             
    .in_ready          (din_ready_0_27),             
    .out_data          (back_data_0_27),              
    .out_valid         (back_valid_0_27),             
    .out_ready         (back_ready_0_27),             
    .fill_level        (din_csr_readdata_0_27),
    .almost_full       (din_almost_full_0_27),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_28"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_28 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_28_r2),              
    .in_valid          (din_valid_0_28_r2),             
    .in_ready          (din_ready_0_28),             
    .out_data          (back_data_0_28),              
    .out_valid         (back_valid_0_28),             
    .out_ready         (back_ready_0_28),             
    .fill_level        (din_csr_readdata_0_28),
    .almost_full       (din_almost_full_0_28),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_29"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_29 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_29_r2),              
    .in_valid          (din_valid_0_29_r2),             
    .in_ready          (din_ready_0_29),             
    .out_data          (back_data_0_29),              
    .out_valid         (back_valid_0_29),             
    .out_ready         (back_ready_0_29),             
    .fill_level        (din_csr_readdata_0_29),
    .almost_full       (din_almost_full_0_29),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_30"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_30 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_30_r2),              
    .in_valid          (din_valid_0_30_r2),             
    .in_ready          (din_ready_0_30),             
    .out_data          (back_data_0_30),              
    .out_valid         (back_valid_0_30),             
    .out_ready         (back_ready_0_30),             
    .fill_level        (din_csr_readdata_0_30),
    .almost_full       (din_almost_full_0_30),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_0_31"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_0_31 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_0_31_r2),              
    .in_valid          (din_valid_0_31_r2),             
    .in_ready          (din_ready_0_31),             
    .out_data          (back_data_0_31),              
    .out_valid         (back_valid_0_31),             
    .out_ready         (back_ready_0_31),             
    .fill_level        (din_csr_readdata_0_31),
    .almost_full       (din_almost_full_0_31),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_0"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_0 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_0_r2),              
    .in_valid          (din_valid_1_0_r2),             
    .in_ready          (din_ready_1_0),             
    .out_data          (back_data_1_0),              
    .out_valid         (back_valid_1_0),             
    .out_ready         (back_ready_1_0),             
    .fill_level        (din_csr_readdata_1_0),
    .almost_full       (din_almost_full_1_0),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_1"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_1 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_1_r2),              
    .in_valid          (din_valid_1_1_r2),             
    .in_ready          (din_ready_1_1),             
    .out_data          (back_data_1_1),              
    .out_valid         (back_valid_1_1),             
    .out_ready         (back_ready_1_1),             
    .fill_level        (din_csr_readdata_1_1),
    .almost_full       (din_almost_full_1_1),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_2"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_2 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_2_r2),              
    .in_valid          (din_valid_1_2_r2),             
    .in_ready          (din_ready_1_2),             
    .out_data          (back_data_1_2),              
    .out_valid         (back_valid_1_2),             
    .out_ready         (back_ready_1_2),             
    .fill_level        (din_csr_readdata_1_2),
    .almost_full       (din_almost_full_1_2),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_3"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_3 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_3_r2),              
    .in_valid          (din_valid_1_3_r2),             
    .in_ready          (din_ready_1_3),             
    .out_data          (back_data_1_3),              
    .out_valid         (back_valid_1_3),             
    .out_ready         (back_ready_1_3),             
    .fill_level        (din_csr_readdata_1_3),
    .almost_full       (din_almost_full_1_3),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_4"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_4 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_4_r2),              
    .in_valid          (din_valid_1_4_r2),             
    .in_ready          (din_ready_1_4),             
    .out_data          (back_data_1_4),              
    .out_valid         (back_valid_1_4),             
    .out_ready         (back_ready_1_4),             
    .fill_level        (din_csr_readdata_1_4),
    .almost_full       (din_almost_full_1_4),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_5"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_5 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_5_r2),              
    .in_valid          (din_valid_1_5_r2),             
    .in_ready          (din_ready_1_5),             
    .out_data          (back_data_1_5),              
    .out_valid         (back_valid_1_5),             
    .out_ready         (back_ready_1_5),             
    .fill_level        (din_csr_readdata_1_5),
    .almost_full       (din_almost_full_1_5),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_6"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_6 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_6_r2),              
    .in_valid          (din_valid_1_6_r2),             
    .in_ready          (din_ready_1_6),             
    .out_data          (back_data_1_6),              
    .out_valid         (back_valid_1_6),             
    .out_ready         (back_ready_1_6),             
    .fill_level        (din_csr_readdata_1_6),
    .almost_full       (din_almost_full_1_6),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_7"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_7 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_7_r2),              
    .in_valid          (din_valid_1_7_r2),             
    .in_ready          (din_ready_1_7),             
    .out_data          (back_data_1_7),              
    .out_valid         (back_valid_1_7),             
    .out_ready         (back_ready_1_7),             
    .fill_level        (din_csr_readdata_1_7),
    .almost_full       (din_almost_full_1_7),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_8"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_8 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_8_r2),              
    .in_valid          (din_valid_1_8_r2),             
    .in_ready          (din_ready_1_8),             
    .out_data          (back_data_1_8),              
    .out_valid         (back_valid_1_8),             
    .out_ready         (back_ready_1_8),             
    .fill_level        (din_csr_readdata_1_8),
    .almost_full       (din_almost_full_1_8),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_9"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_9 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_9_r2),              
    .in_valid          (din_valid_1_9_r2),             
    .in_ready          (din_ready_1_9),             
    .out_data          (back_data_1_9),              
    .out_valid         (back_valid_1_9),             
    .out_ready         (back_ready_1_9),             
    .fill_level        (din_csr_readdata_1_9),
    .almost_full       (din_almost_full_1_9),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_10"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_10 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_10_r2),              
    .in_valid          (din_valid_1_10_r2),             
    .in_ready          (din_ready_1_10),             
    .out_data          (back_data_1_10),              
    .out_valid         (back_valid_1_10),             
    .out_ready         (back_ready_1_10),             
    .fill_level        (din_csr_readdata_1_10),
    .almost_full       (din_almost_full_1_10),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_11"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_11 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_11_r2),              
    .in_valid          (din_valid_1_11_r2),             
    .in_ready          (din_ready_1_11),             
    .out_data          (back_data_1_11),              
    .out_valid         (back_valid_1_11),             
    .out_ready         (back_ready_1_11),             
    .fill_level        (din_csr_readdata_1_11),
    .almost_full       (din_almost_full_1_11),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_12"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_12 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_12_r2),              
    .in_valid          (din_valid_1_12_r2),             
    .in_ready          (din_ready_1_12),             
    .out_data          (back_data_1_12),              
    .out_valid         (back_valid_1_12),             
    .out_ready         (back_ready_1_12),             
    .fill_level        (din_csr_readdata_1_12),
    .almost_full       (din_almost_full_1_12),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_13"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_13 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_13_r2),              
    .in_valid          (din_valid_1_13_r2),             
    .in_ready          (din_ready_1_13),             
    .out_data          (back_data_1_13),              
    .out_valid         (back_valid_1_13),             
    .out_ready         (back_ready_1_13),             
    .fill_level        (din_csr_readdata_1_13),
    .almost_full       (din_almost_full_1_13),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_14"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_14 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_14_r2),              
    .in_valid          (din_valid_1_14_r2),             
    .in_ready          (din_ready_1_14),             
    .out_data          (back_data_1_14),              
    .out_valid         (back_valid_1_14),             
    .out_ready         (back_ready_1_14),             
    .fill_level        (din_csr_readdata_1_14),
    .almost_full       (din_almost_full_1_14),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_15"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_15 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_15_r2),              
    .in_valid          (din_valid_1_15_r2),             
    .in_ready          (din_ready_1_15),             
    .out_data          (back_data_1_15),              
    .out_valid         (back_valid_1_15),             
    .out_ready         (back_ready_1_15),             
    .fill_level        (din_csr_readdata_1_15),
    .almost_full       (din_almost_full_1_15),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_16"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_16 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_16_r2),              
    .in_valid          (din_valid_1_16_r2),             
    .in_ready          (din_ready_1_16),             
    .out_data          (back_data_1_16),              
    .out_valid         (back_valid_1_16),             
    .out_ready         (back_ready_1_16),             
    .fill_level        (din_csr_readdata_1_16),
    .almost_full       (din_almost_full_1_16),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_17"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_17 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_17_r2),              
    .in_valid          (din_valid_1_17_r2),             
    .in_ready          (din_ready_1_17),             
    .out_data          (back_data_1_17),              
    .out_valid         (back_valid_1_17),             
    .out_ready         (back_ready_1_17),             
    .fill_level        (din_csr_readdata_1_17),
    .almost_full       (din_almost_full_1_17),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_18"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_18 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_18_r2),              
    .in_valid          (din_valid_1_18_r2),             
    .in_ready          (din_ready_1_18),             
    .out_data          (back_data_1_18),              
    .out_valid         (back_valid_1_18),             
    .out_ready         (back_ready_1_18),             
    .fill_level        (din_csr_readdata_1_18),
    .almost_full       (din_almost_full_1_18),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_19"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_19 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_19_r2),              
    .in_valid          (din_valid_1_19_r2),             
    .in_ready          (din_ready_1_19),             
    .out_data          (back_data_1_19),              
    .out_valid         (back_valid_1_19),             
    .out_ready         (back_ready_1_19),             
    .fill_level        (din_csr_readdata_1_19),
    .almost_full       (din_almost_full_1_19),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_20"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_20 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_20_r2),              
    .in_valid          (din_valid_1_20_r2),             
    .in_ready          (din_ready_1_20),             
    .out_data          (back_data_1_20),              
    .out_valid         (back_valid_1_20),             
    .out_ready         (back_ready_1_20),             
    .fill_level        (din_csr_readdata_1_20),
    .almost_full       (din_almost_full_1_20),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_21"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_21 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_21_r2),              
    .in_valid          (din_valid_1_21_r2),             
    .in_ready          (din_ready_1_21),             
    .out_data          (back_data_1_21),              
    .out_valid         (back_valid_1_21),             
    .out_ready         (back_ready_1_21),             
    .fill_level        (din_csr_readdata_1_21),
    .almost_full       (din_almost_full_1_21),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_22"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_22 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_22_r2),              
    .in_valid          (din_valid_1_22_r2),             
    .in_ready          (din_ready_1_22),             
    .out_data          (back_data_1_22),              
    .out_valid         (back_valid_1_22),             
    .out_ready         (back_ready_1_22),             
    .fill_level        (din_csr_readdata_1_22),
    .almost_full       (din_almost_full_1_22),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_23"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_23 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_23_r2),              
    .in_valid          (din_valid_1_23_r2),             
    .in_ready          (din_ready_1_23),             
    .out_data          (back_data_1_23),              
    .out_valid         (back_valid_1_23),             
    .out_ready         (back_ready_1_23),             
    .fill_level        (din_csr_readdata_1_23),
    .almost_full       (din_almost_full_1_23),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_24"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_24 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_24_r2),              
    .in_valid          (din_valid_1_24_r2),             
    .in_ready          (din_ready_1_24),             
    .out_data          (back_data_1_24),              
    .out_valid         (back_valid_1_24),             
    .out_ready         (back_ready_1_24),             
    .fill_level        (din_csr_readdata_1_24),
    .almost_full       (din_almost_full_1_24),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_25"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_25 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_25_r2),              
    .in_valid          (din_valid_1_25_r2),             
    .in_ready          (din_ready_1_25),             
    .out_data          (back_data_1_25),              
    .out_valid         (back_valid_1_25),             
    .out_ready         (back_ready_1_25),             
    .fill_level        (din_csr_readdata_1_25),
    .almost_full       (din_almost_full_1_25),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_26"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_26 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_26_r2),              
    .in_valid          (din_valid_1_26_r2),             
    .in_ready          (din_ready_1_26),             
    .out_data          (back_data_1_26),              
    .out_valid         (back_valid_1_26),             
    .out_ready         (back_ready_1_26),             
    .fill_level        (din_csr_readdata_1_26),
    .almost_full       (din_almost_full_1_26),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_27"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_27 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_27_r2),              
    .in_valid          (din_valid_1_27_r2),             
    .in_ready          (din_ready_1_27),             
    .out_data          (back_data_1_27),              
    .out_valid         (back_valid_1_27),             
    .out_ready         (back_ready_1_27),             
    .fill_level        (din_csr_readdata_1_27),
    .almost_full       (din_almost_full_1_27),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_28"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_28 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_28_r2),              
    .in_valid          (din_valid_1_28_r2),             
    .in_ready          (din_ready_1_28),             
    .out_data          (back_data_1_28),              
    .out_valid         (back_valid_1_28),             
    .out_ready         (back_ready_1_28),             
    .fill_level        (din_csr_readdata_1_28),
    .almost_full       (din_almost_full_1_28),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_29"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_29 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_29_r2),              
    .in_valid          (din_valid_1_29_r2),             
    .in_ready          (din_ready_1_29),             
    .out_data          (back_data_1_29),              
    .out_valid         (back_valid_1_29),             
    .out_ready         (back_ready_1_29),             
    .fill_level        (din_csr_readdata_1_29),
    .almost_full       (din_almost_full_1_29),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_30"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_30 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_30_r2),              
    .in_valid          (din_valid_1_30_r2),             
    .in_ready          (din_ready_1_30),             
    .out_data          (back_data_1_30),              
    .out_valid         (back_valid_1_30),             
    .out_ready         (back_ready_1_30),             
    .fill_level        (din_csr_readdata_1_30),
    .almost_full       (din_almost_full_1_30),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_1_31"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_1_31 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_1_31_r2),              
    .in_valid          (din_valid_1_31_r2),             
    .in_ready          (din_ready_1_31),             
    .out_data          (back_data_1_31),              
    .out_valid         (back_valid_1_31),             
    .out_ready         (back_ready_1_31),             
    .fill_level        (din_csr_readdata_1_31),
    .almost_full       (din_almost_full_1_31),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_0"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_0 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_0_r2),              
    .in_valid          (din_valid_2_0_r2),             
    .in_ready          (din_ready_2_0),             
    .out_data          (back_data_2_0),              
    .out_valid         (back_valid_2_0),             
    .out_ready         (back_ready_2_0),             
    .fill_level        (din_csr_readdata_2_0),
    .almost_full       (din_almost_full_2_0),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_1"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_1 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_1_r2),              
    .in_valid          (din_valid_2_1_r2),             
    .in_ready          (din_ready_2_1),             
    .out_data          (back_data_2_1),              
    .out_valid         (back_valid_2_1),             
    .out_ready         (back_ready_2_1),             
    .fill_level        (din_csr_readdata_2_1),
    .almost_full       (din_almost_full_2_1),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_2"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_2 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_2_r2),              
    .in_valid          (din_valid_2_2_r2),             
    .in_ready          (din_ready_2_2),             
    .out_data          (back_data_2_2),              
    .out_valid         (back_valid_2_2),             
    .out_ready         (back_ready_2_2),             
    .fill_level        (din_csr_readdata_2_2),
    .almost_full       (din_almost_full_2_2),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_3"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_3 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_3_r2),              
    .in_valid          (din_valid_2_3_r2),             
    .in_ready          (din_ready_2_3),             
    .out_data          (back_data_2_3),              
    .out_valid         (back_valid_2_3),             
    .out_ready         (back_ready_2_3),             
    .fill_level        (din_csr_readdata_2_3),
    .almost_full       (din_almost_full_2_3),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_4"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_4 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_4_r2),              
    .in_valid          (din_valid_2_4_r2),             
    .in_ready          (din_ready_2_4),             
    .out_data          (back_data_2_4),              
    .out_valid         (back_valid_2_4),             
    .out_ready         (back_ready_2_4),             
    .fill_level        (din_csr_readdata_2_4),
    .almost_full       (din_almost_full_2_4),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_5"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_5 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_5_r2),              
    .in_valid          (din_valid_2_5_r2),             
    .in_ready          (din_ready_2_5),             
    .out_data          (back_data_2_5),              
    .out_valid         (back_valid_2_5),             
    .out_ready         (back_ready_2_5),             
    .fill_level        (din_csr_readdata_2_5),
    .almost_full       (din_almost_full_2_5),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_6"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_6 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_6_r2),              
    .in_valid          (din_valid_2_6_r2),             
    .in_ready          (din_ready_2_6),             
    .out_data          (back_data_2_6),              
    .out_valid         (back_valid_2_6),             
    .out_ready         (back_ready_2_6),             
    .fill_level        (din_csr_readdata_2_6),
    .almost_full       (din_almost_full_2_6),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_7"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_7 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_7_r2),              
    .in_valid          (din_valid_2_7_r2),             
    .in_ready          (din_ready_2_7),             
    .out_data          (back_data_2_7),              
    .out_valid         (back_valid_2_7),             
    .out_ready         (back_ready_2_7),             
    .fill_level        (din_csr_readdata_2_7),
    .almost_full       (din_almost_full_2_7),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_8"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_8 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_8_r2),              
    .in_valid          (din_valid_2_8_r2),             
    .in_ready          (din_ready_2_8),             
    .out_data          (back_data_2_8),              
    .out_valid         (back_valid_2_8),             
    .out_ready         (back_ready_2_8),             
    .fill_level        (din_csr_readdata_2_8),
    .almost_full       (din_almost_full_2_8),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_9"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_9 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_9_r2),              
    .in_valid          (din_valid_2_9_r2),             
    .in_ready          (din_ready_2_9),             
    .out_data          (back_data_2_9),              
    .out_valid         (back_valid_2_9),             
    .out_ready         (back_ready_2_9),             
    .fill_level        (din_csr_readdata_2_9),
    .almost_full       (din_almost_full_2_9),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_10"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_10 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_10_r2),              
    .in_valid          (din_valid_2_10_r2),             
    .in_ready          (din_ready_2_10),             
    .out_data          (back_data_2_10),              
    .out_valid         (back_valid_2_10),             
    .out_ready         (back_ready_2_10),             
    .fill_level        (din_csr_readdata_2_10),
    .almost_full       (din_almost_full_2_10),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_11"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_11 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_11_r2),              
    .in_valid          (din_valid_2_11_r2),             
    .in_ready          (din_ready_2_11),             
    .out_data          (back_data_2_11),              
    .out_valid         (back_valid_2_11),             
    .out_ready         (back_ready_2_11),             
    .fill_level        (din_csr_readdata_2_11),
    .almost_full       (din_almost_full_2_11),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_12"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_12 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_12_r2),              
    .in_valid          (din_valid_2_12_r2),             
    .in_ready          (din_ready_2_12),             
    .out_data          (back_data_2_12),              
    .out_valid         (back_valid_2_12),             
    .out_ready         (back_ready_2_12),             
    .fill_level        (din_csr_readdata_2_12),
    .almost_full       (din_almost_full_2_12),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_13"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_13 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_13_r2),              
    .in_valid          (din_valid_2_13_r2),             
    .in_ready          (din_ready_2_13),             
    .out_data          (back_data_2_13),              
    .out_valid         (back_valid_2_13),             
    .out_ready         (back_ready_2_13),             
    .fill_level        (din_csr_readdata_2_13),
    .almost_full       (din_almost_full_2_13),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_14"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_14 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_14_r2),              
    .in_valid          (din_valid_2_14_r2),             
    .in_ready          (din_ready_2_14),             
    .out_data          (back_data_2_14),              
    .out_valid         (back_valid_2_14),             
    .out_ready         (back_ready_2_14),             
    .fill_level        (din_csr_readdata_2_14),
    .almost_full       (din_almost_full_2_14),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_15"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_15 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_15_r2),              
    .in_valid          (din_valid_2_15_r2),             
    .in_ready          (din_ready_2_15),             
    .out_data          (back_data_2_15),              
    .out_valid         (back_valid_2_15),             
    .out_ready         (back_ready_2_15),             
    .fill_level        (din_csr_readdata_2_15),
    .almost_full       (din_almost_full_2_15),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_16"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_16 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_16_r2),              
    .in_valid          (din_valid_2_16_r2),             
    .in_ready          (din_ready_2_16),             
    .out_data          (back_data_2_16),              
    .out_valid         (back_valid_2_16),             
    .out_ready         (back_ready_2_16),             
    .fill_level        (din_csr_readdata_2_16),
    .almost_full       (din_almost_full_2_16),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_17"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_17 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_17_r2),              
    .in_valid          (din_valid_2_17_r2),             
    .in_ready          (din_ready_2_17),             
    .out_data          (back_data_2_17),              
    .out_valid         (back_valid_2_17),             
    .out_ready         (back_ready_2_17),             
    .fill_level        (din_csr_readdata_2_17),
    .almost_full       (din_almost_full_2_17),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_18"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_18 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_18_r2),              
    .in_valid          (din_valid_2_18_r2),             
    .in_ready          (din_ready_2_18),             
    .out_data          (back_data_2_18),              
    .out_valid         (back_valid_2_18),             
    .out_ready         (back_ready_2_18),             
    .fill_level        (din_csr_readdata_2_18),
    .almost_full       (din_almost_full_2_18),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_19"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_19 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_19_r2),              
    .in_valid          (din_valid_2_19_r2),             
    .in_ready          (din_ready_2_19),             
    .out_data          (back_data_2_19),              
    .out_valid         (back_valid_2_19),             
    .out_ready         (back_ready_2_19),             
    .fill_level        (din_csr_readdata_2_19),
    .almost_full       (din_almost_full_2_19),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_20"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_20 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_20_r2),              
    .in_valid          (din_valid_2_20_r2),             
    .in_ready          (din_ready_2_20),             
    .out_data          (back_data_2_20),              
    .out_valid         (back_valid_2_20),             
    .out_ready         (back_ready_2_20),             
    .fill_level        (din_csr_readdata_2_20),
    .almost_full       (din_almost_full_2_20),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_21"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_21 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_21_r2),              
    .in_valid          (din_valid_2_21_r2),             
    .in_ready          (din_ready_2_21),             
    .out_data          (back_data_2_21),              
    .out_valid         (back_valid_2_21),             
    .out_ready         (back_ready_2_21),             
    .fill_level        (din_csr_readdata_2_21),
    .almost_full       (din_almost_full_2_21),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_22"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_22 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_22_r2),              
    .in_valid          (din_valid_2_22_r2),             
    .in_ready          (din_ready_2_22),             
    .out_data          (back_data_2_22),              
    .out_valid         (back_valid_2_22),             
    .out_ready         (back_ready_2_22),             
    .fill_level        (din_csr_readdata_2_22),
    .almost_full       (din_almost_full_2_22),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_23"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_23 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_23_r2),              
    .in_valid          (din_valid_2_23_r2),             
    .in_ready          (din_ready_2_23),             
    .out_data          (back_data_2_23),              
    .out_valid         (back_valid_2_23),             
    .out_ready         (back_ready_2_23),             
    .fill_level        (din_csr_readdata_2_23),
    .almost_full       (din_almost_full_2_23),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_24"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_24 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_24_r2),              
    .in_valid          (din_valid_2_24_r2),             
    .in_ready          (din_ready_2_24),             
    .out_data          (back_data_2_24),              
    .out_valid         (back_valid_2_24),             
    .out_ready         (back_ready_2_24),             
    .fill_level        (din_csr_readdata_2_24),
    .almost_full       (din_almost_full_2_24),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_25"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_25 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_25_r2),              
    .in_valid          (din_valid_2_25_r2),             
    .in_ready          (din_ready_2_25),             
    .out_data          (back_data_2_25),              
    .out_valid         (back_valid_2_25),             
    .out_ready         (back_ready_2_25),             
    .fill_level        (din_csr_readdata_2_25),
    .almost_full       (din_almost_full_2_25),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_26"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_26 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_26_r2),              
    .in_valid          (din_valid_2_26_r2),             
    .in_ready          (din_ready_2_26),             
    .out_data          (back_data_2_26),              
    .out_valid         (back_valid_2_26),             
    .out_ready         (back_ready_2_26),             
    .fill_level        (din_csr_readdata_2_26),
    .almost_full       (din_almost_full_2_26),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_27"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_27 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_27_r2),              
    .in_valid          (din_valid_2_27_r2),             
    .in_ready          (din_ready_2_27),             
    .out_data          (back_data_2_27),              
    .out_valid         (back_valid_2_27),             
    .out_ready         (back_ready_2_27),             
    .fill_level        (din_csr_readdata_2_27),
    .almost_full       (din_almost_full_2_27),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_28"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_28 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_28_r2),              
    .in_valid          (din_valid_2_28_r2),             
    .in_ready          (din_ready_2_28),             
    .out_data          (back_data_2_28),              
    .out_valid         (back_valid_2_28),             
    .out_ready         (back_ready_2_28),             
    .fill_level        (din_csr_readdata_2_28),
    .almost_full       (din_almost_full_2_28),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_29"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_29 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_29_r2),              
    .in_valid          (din_valid_2_29_r2),             
    .in_ready          (din_ready_2_29),             
    .out_data          (back_data_2_29),              
    .out_valid         (back_valid_2_29),             
    .out_ready         (back_ready_2_29),             
    .fill_level        (din_csr_readdata_2_29),
    .almost_full       (din_almost_full_2_29),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_30"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_30 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_30_r2),              
    .in_valid          (din_valid_2_30_r2),             
    .in_ready          (din_ready_2_30),             
    .out_data          (back_data_2_30),              
    .out_valid         (back_valid_2_30),             
    .out_ready         (back_ready_2_30),             
    .fill_level        (din_csr_readdata_2_30),
    .almost_full       (din_almost_full_2_30),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_2_31"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_2_31 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_2_31_r2),              
    .in_valid          (din_valid_2_31_r2),             
    .in_ready          (din_ready_2_31),             
    .out_data          (back_data_2_31),              
    .out_valid         (back_valid_2_31),             
    .out_ready         (back_ready_2_31),             
    .fill_level        (din_csr_readdata_2_31),
    .almost_full       (din_almost_full_2_31),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_0"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_0 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_0_r2),              
    .in_valid          (din_valid_3_0_r2),             
    .in_ready          (din_ready_3_0),             
    .out_data          (back_data_3_0),              
    .out_valid         (back_valid_3_0),             
    .out_ready         (back_ready_3_0),             
    .fill_level        (din_csr_readdata_3_0),
    .almost_full       (din_almost_full_3_0),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_1"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_1 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_1_r2),              
    .in_valid          (din_valid_3_1_r2),             
    .in_ready          (din_ready_3_1),             
    .out_data          (back_data_3_1),              
    .out_valid         (back_valid_3_1),             
    .out_ready         (back_ready_3_1),             
    .fill_level        (din_csr_readdata_3_1),
    .almost_full       (din_almost_full_3_1),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_2"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_2 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_2_r2),              
    .in_valid          (din_valid_3_2_r2),             
    .in_ready          (din_ready_3_2),             
    .out_data          (back_data_3_2),              
    .out_valid         (back_valid_3_2),             
    .out_ready         (back_ready_3_2),             
    .fill_level        (din_csr_readdata_3_2),
    .almost_full       (din_almost_full_3_2),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_3"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_3 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_3_r2),              
    .in_valid          (din_valid_3_3_r2),             
    .in_ready          (din_ready_3_3),             
    .out_data          (back_data_3_3),              
    .out_valid         (back_valid_3_3),             
    .out_ready         (back_ready_3_3),             
    .fill_level        (din_csr_readdata_3_3),
    .almost_full       (din_almost_full_3_3),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_4"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_4 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_4_r2),              
    .in_valid          (din_valid_3_4_r2),             
    .in_ready          (din_ready_3_4),             
    .out_data          (back_data_3_4),              
    .out_valid         (back_valid_3_4),             
    .out_ready         (back_ready_3_4),             
    .fill_level        (din_csr_readdata_3_4),
    .almost_full       (din_almost_full_3_4),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_5"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_5 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_5_r2),              
    .in_valid          (din_valid_3_5_r2),             
    .in_ready          (din_ready_3_5),             
    .out_data          (back_data_3_5),              
    .out_valid         (back_valid_3_5),             
    .out_ready         (back_ready_3_5),             
    .fill_level        (din_csr_readdata_3_5),
    .almost_full       (din_almost_full_3_5),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_6"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_6 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_6_r2),              
    .in_valid          (din_valid_3_6_r2),             
    .in_ready          (din_ready_3_6),             
    .out_data          (back_data_3_6),              
    .out_valid         (back_valid_3_6),             
    .out_ready         (back_ready_3_6),             
    .fill_level        (din_csr_readdata_3_6),
    .almost_full       (din_almost_full_3_6),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_7"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_7 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_7_r2),              
    .in_valid          (din_valid_3_7_r2),             
    .in_ready          (din_ready_3_7),             
    .out_data          (back_data_3_7),              
    .out_valid         (back_valid_3_7),             
    .out_ready         (back_ready_3_7),             
    .fill_level        (din_csr_readdata_3_7),
    .almost_full       (din_almost_full_3_7),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_8"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_8 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_8_r2),              
    .in_valid          (din_valid_3_8_r2),             
    .in_ready          (din_ready_3_8),             
    .out_data          (back_data_3_8),              
    .out_valid         (back_valid_3_8),             
    .out_ready         (back_ready_3_8),             
    .fill_level        (din_csr_readdata_3_8),
    .almost_full       (din_almost_full_3_8),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_9"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_9 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_9_r2),              
    .in_valid          (din_valid_3_9_r2),             
    .in_ready          (din_ready_3_9),             
    .out_data          (back_data_3_9),              
    .out_valid         (back_valid_3_9),             
    .out_ready         (back_ready_3_9),             
    .fill_level        (din_csr_readdata_3_9),
    .almost_full       (din_almost_full_3_9),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_10"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_10 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_10_r2),              
    .in_valid          (din_valid_3_10_r2),             
    .in_ready          (din_ready_3_10),             
    .out_data          (back_data_3_10),              
    .out_valid         (back_valid_3_10),             
    .out_ready         (back_ready_3_10),             
    .fill_level        (din_csr_readdata_3_10),
    .almost_full       (din_almost_full_3_10),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_11"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_11 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_11_r2),              
    .in_valid          (din_valid_3_11_r2),             
    .in_ready          (din_ready_3_11),             
    .out_data          (back_data_3_11),              
    .out_valid         (back_valid_3_11),             
    .out_ready         (back_ready_3_11),             
    .fill_level        (din_csr_readdata_3_11),
    .almost_full       (din_almost_full_3_11),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_12"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_12 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_12_r2),              
    .in_valid          (din_valid_3_12_r2),             
    .in_ready          (din_ready_3_12),             
    .out_data          (back_data_3_12),              
    .out_valid         (back_valid_3_12),             
    .out_ready         (back_ready_3_12),             
    .fill_level        (din_csr_readdata_3_12),
    .almost_full       (din_almost_full_3_12),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_13"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_13 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_13_r2),              
    .in_valid          (din_valid_3_13_r2),             
    .in_ready          (din_ready_3_13),             
    .out_data          (back_data_3_13),              
    .out_valid         (back_valid_3_13),             
    .out_ready         (back_ready_3_13),             
    .fill_level        (din_csr_readdata_3_13),
    .almost_full       (din_almost_full_3_13),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_14"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_14 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_14_r2),              
    .in_valid          (din_valid_3_14_r2),             
    .in_ready          (din_ready_3_14),             
    .out_data          (back_data_3_14),              
    .out_valid         (back_valid_3_14),             
    .out_ready         (back_ready_3_14),             
    .fill_level        (din_csr_readdata_3_14),
    .almost_full       (din_almost_full_3_14),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_15"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_15 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_15_r2),              
    .in_valid          (din_valid_3_15_r2),             
    .in_ready          (din_ready_3_15),             
    .out_data          (back_data_3_15),              
    .out_valid         (back_valid_3_15),             
    .out_ready         (back_ready_3_15),             
    .fill_level        (din_csr_readdata_3_15),
    .almost_full       (din_almost_full_3_15),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_16"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_16 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_16_r2),              
    .in_valid          (din_valid_3_16_r2),             
    .in_ready          (din_ready_3_16),             
    .out_data          (back_data_3_16),              
    .out_valid         (back_valid_3_16),             
    .out_ready         (back_ready_3_16),             
    .fill_level        (din_csr_readdata_3_16),
    .almost_full       (din_almost_full_3_16),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_17"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_17 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_17_r2),              
    .in_valid          (din_valid_3_17_r2),             
    .in_ready          (din_ready_3_17),             
    .out_data          (back_data_3_17),              
    .out_valid         (back_valid_3_17),             
    .out_ready         (back_ready_3_17),             
    .fill_level        (din_csr_readdata_3_17),
    .almost_full       (din_almost_full_3_17),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_18"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_18 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_18_r2),              
    .in_valid          (din_valid_3_18_r2),             
    .in_ready          (din_ready_3_18),             
    .out_data          (back_data_3_18),              
    .out_valid         (back_valid_3_18),             
    .out_ready         (back_ready_3_18),             
    .fill_level        (din_csr_readdata_3_18),
    .almost_full       (din_almost_full_3_18),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_19"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_19 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_19_r2),              
    .in_valid          (din_valid_3_19_r2),             
    .in_ready          (din_ready_3_19),             
    .out_data          (back_data_3_19),              
    .out_valid         (back_valid_3_19),             
    .out_ready         (back_ready_3_19),             
    .fill_level        (din_csr_readdata_3_19),
    .almost_full       (din_almost_full_3_19),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_20"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_20 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_20_r2),              
    .in_valid          (din_valid_3_20_r2),             
    .in_ready          (din_ready_3_20),             
    .out_data          (back_data_3_20),              
    .out_valid         (back_valid_3_20),             
    .out_ready         (back_ready_3_20),             
    .fill_level        (din_csr_readdata_3_20),
    .almost_full       (din_almost_full_3_20),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_21"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_21 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_21_r2),              
    .in_valid          (din_valid_3_21_r2),             
    .in_ready          (din_ready_3_21),             
    .out_data          (back_data_3_21),              
    .out_valid         (back_valid_3_21),             
    .out_ready         (back_ready_3_21),             
    .fill_level        (din_csr_readdata_3_21),
    .almost_full       (din_almost_full_3_21),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_22"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_22 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_22_r2),              
    .in_valid          (din_valid_3_22_r2),             
    .in_ready          (din_ready_3_22),             
    .out_data          (back_data_3_22),              
    .out_valid         (back_valid_3_22),             
    .out_ready         (back_ready_3_22),             
    .fill_level        (din_csr_readdata_3_22),
    .almost_full       (din_almost_full_3_22),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_23"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_23 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_23_r2),              
    .in_valid          (din_valid_3_23_r2),             
    .in_ready          (din_ready_3_23),             
    .out_data          (back_data_3_23),              
    .out_valid         (back_valid_3_23),             
    .out_ready         (back_ready_3_23),             
    .fill_level        (din_csr_readdata_3_23),
    .almost_full       (din_almost_full_3_23),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_24"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_24 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_24_r2),              
    .in_valid          (din_valid_3_24_r2),             
    .in_ready          (din_ready_3_24),             
    .out_data          (back_data_3_24),              
    .out_valid         (back_valid_3_24),             
    .out_ready         (back_ready_3_24),             
    .fill_level        (din_csr_readdata_3_24),
    .almost_full       (din_almost_full_3_24),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_25"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_25 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_25_r2),              
    .in_valid          (din_valid_3_25_r2),             
    .in_ready          (din_ready_3_25),             
    .out_data          (back_data_3_25),              
    .out_valid         (back_valid_3_25),             
    .out_ready         (back_ready_3_25),             
    .fill_level        (din_csr_readdata_3_25),
    .almost_full       (din_almost_full_3_25),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_26"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_26 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_26_r2),              
    .in_valid          (din_valid_3_26_r2),             
    .in_ready          (din_ready_3_26),             
    .out_data          (back_data_3_26),              
    .out_valid         (back_valid_3_26),             
    .out_ready         (back_ready_3_26),             
    .fill_level        (din_csr_readdata_3_26),
    .almost_full       (din_almost_full_3_26),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_27"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_27 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_27_r2),              
    .in_valid          (din_valid_3_27_r2),             
    .in_ready          (din_ready_3_27),             
    .out_data          (back_data_3_27),              
    .out_valid         (back_valid_3_27),             
    .out_ready         (back_ready_3_27),             
    .fill_level        (din_csr_readdata_3_27),
    .almost_full       (din_almost_full_3_27),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_28"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_28 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_28_r2),              
    .in_valid          (din_valid_3_28_r2),             
    .in_ready          (din_ready_3_28),             
    .out_data          (back_data_3_28),              
    .out_valid         (back_valid_3_28),             
    .out_ready         (back_ready_3_28),             
    .fill_level        (din_csr_readdata_3_28),
    .almost_full       (din_almost_full_3_28),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_29"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_29 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_29_r2),              
    .in_valid          (din_valid_3_29_r2),             
    .in_ready          (din_ready_3_29),             
    .out_data          (back_data_3_29),              
    .out_valid         (back_valid_3_29),             
    .out_ready         (back_ready_3_29),             
    .fill_level        (din_csr_readdata_3_29),
    .almost_full       (din_almost_full_3_29),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_30"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_30 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_30_r2),              
    .in_valid          (din_valid_3_30_r2),             
    .in_ready          (din_ready_3_30),             
    .out_data          (back_data_3_30),              
    .out_valid         (back_valid_3_30),             
    .out_ready         (back_ready_3_30),             
    .fill_level        (din_csr_readdata_3_30),
    .almost_full       (din_almost_full_3_30),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_3_31"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_3_31 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_3_31_r2),              
    .in_valid          (din_valid_3_31_r2),             
    .in_ready          (din_ready_3_31),             
    .out_data          (back_data_3_31),              
    .out_valid         (back_valid_3_31),             
    .out_ready         (back_ready_3_31),             
    .fill_level        (din_csr_readdata_3_31),
    .almost_full       (din_almost_full_3_31),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_0"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_0 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_0_r2),              
    .in_valid          (din_valid_4_0_r2),             
    .in_ready          (din_ready_4_0),             
    .out_data          (back_data_4_0),              
    .out_valid         (back_valid_4_0),             
    .out_ready         (back_ready_4_0),             
    .fill_level        (din_csr_readdata_4_0),
    .almost_full       (din_almost_full_4_0),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_1"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_1 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_1_r2),              
    .in_valid          (din_valid_4_1_r2),             
    .in_ready          (din_ready_4_1),             
    .out_data          (back_data_4_1),              
    .out_valid         (back_valid_4_1),             
    .out_ready         (back_ready_4_1),             
    .fill_level        (din_csr_readdata_4_1),
    .almost_full       (din_almost_full_4_1),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_2"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_2 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_2_r2),              
    .in_valid          (din_valid_4_2_r2),             
    .in_ready          (din_ready_4_2),             
    .out_data          (back_data_4_2),              
    .out_valid         (back_valid_4_2),             
    .out_ready         (back_ready_4_2),             
    .fill_level        (din_csr_readdata_4_2),
    .almost_full       (din_almost_full_4_2),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_3"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_3 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_3_r2),              
    .in_valid          (din_valid_4_3_r2),             
    .in_ready          (din_ready_4_3),             
    .out_data          (back_data_4_3),              
    .out_valid         (back_valid_4_3),             
    .out_ready         (back_ready_4_3),             
    .fill_level        (din_csr_readdata_4_3),
    .almost_full       (din_almost_full_4_3),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_4"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_4 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_4_r2),              
    .in_valid          (din_valid_4_4_r2),             
    .in_ready          (din_ready_4_4),             
    .out_data          (back_data_4_4),              
    .out_valid         (back_valid_4_4),             
    .out_ready         (back_ready_4_4),             
    .fill_level        (din_csr_readdata_4_4),
    .almost_full       (din_almost_full_4_4),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_5"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_5 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_5_r2),              
    .in_valid          (din_valid_4_5_r2),             
    .in_ready          (din_ready_4_5),             
    .out_data          (back_data_4_5),              
    .out_valid         (back_valid_4_5),             
    .out_ready         (back_ready_4_5),             
    .fill_level        (din_csr_readdata_4_5),
    .almost_full       (din_almost_full_4_5),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_6"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_6 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_6_r2),              
    .in_valid          (din_valid_4_6_r2),             
    .in_ready          (din_ready_4_6),             
    .out_data          (back_data_4_6),              
    .out_valid         (back_valid_4_6),             
    .out_ready         (back_ready_4_6),             
    .fill_level        (din_csr_readdata_4_6),
    .almost_full       (din_almost_full_4_6),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_7"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_7 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_7_r2),              
    .in_valid          (din_valid_4_7_r2),             
    .in_ready          (din_ready_4_7),             
    .out_data          (back_data_4_7),              
    .out_valid         (back_valid_4_7),             
    .out_ready         (back_ready_4_7),             
    .fill_level        (din_csr_readdata_4_7),
    .almost_full       (din_almost_full_4_7),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_8"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_8 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_8_r2),              
    .in_valid          (din_valid_4_8_r2),             
    .in_ready          (din_ready_4_8),             
    .out_data          (back_data_4_8),              
    .out_valid         (back_valid_4_8),             
    .out_ready         (back_ready_4_8),             
    .fill_level        (din_csr_readdata_4_8),
    .almost_full       (din_almost_full_4_8),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_9"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_9 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_9_r2),              
    .in_valid          (din_valid_4_9_r2),             
    .in_ready          (din_ready_4_9),             
    .out_data          (back_data_4_9),              
    .out_valid         (back_valid_4_9),             
    .out_ready         (back_ready_4_9),             
    .fill_level        (din_csr_readdata_4_9),
    .almost_full       (din_almost_full_4_9),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_10"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_10 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_10_r2),              
    .in_valid          (din_valid_4_10_r2),             
    .in_ready          (din_ready_4_10),             
    .out_data          (back_data_4_10),              
    .out_valid         (back_valid_4_10),             
    .out_ready         (back_ready_4_10),             
    .fill_level        (din_csr_readdata_4_10),
    .almost_full       (din_almost_full_4_10),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_11"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_11 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_11_r2),              
    .in_valid          (din_valid_4_11_r2),             
    .in_ready          (din_ready_4_11),             
    .out_data          (back_data_4_11),              
    .out_valid         (back_valid_4_11),             
    .out_ready         (back_ready_4_11),             
    .fill_level        (din_csr_readdata_4_11),
    .almost_full       (din_almost_full_4_11),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_12"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_12 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_12_r2),              
    .in_valid          (din_valid_4_12_r2),             
    .in_ready          (din_ready_4_12),             
    .out_data          (back_data_4_12),              
    .out_valid         (back_valid_4_12),             
    .out_ready         (back_ready_4_12),             
    .fill_level        (din_csr_readdata_4_12),
    .almost_full       (din_almost_full_4_12),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_13"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_13 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_13_r2),              
    .in_valid          (din_valid_4_13_r2),             
    .in_ready          (din_ready_4_13),             
    .out_data          (back_data_4_13),              
    .out_valid         (back_valid_4_13),             
    .out_ready         (back_ready_4_13),             
    .fill_level        (din_csr_readdata_4_13),
    .almost_full       (din_almost_full_4_13),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_14"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_14 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_14_r2),              
    .in_valid          (din_valid_4_14_r2),             
    .in_ready          (din_ready_4_14),             
    .out_data          (back_data_4_14),              
    .out_valid         (back_valid_4_14),             
    .out_ready         (back_ready_4_14),             
    .fill_level        (din_csr_readdata_4_14),
    .almost_full       (din_almost_full_4_14),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_15"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_15 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_15_r2),              
    .in_valid          (din_valid_4_15_r2),             
    .in_ready          (din_ready_4_15),             
    .out_data          (back_data_4_15),              
    .out_valid         (back_valid_4_15),             
    .out_ready         (back_ready_4_15),             
    .fill_level        (din_csr_readdata_4_15),
    .almost_full       (din_almost_full_4_15),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_16"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_16 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_16_r2),              
    .in_valid          (din_valid_4_16_r2),             
    .in_ready          (din_ready_4_16),             
    .out_data          (back_data_4_16),              
    .out_valid         (back_valid_4_16),             
    .out_ready         (back_ready_4_16),             
    .fill_level        (din_csr_readdata_4_16),
    .almost_full       (din_almost_full_4_16),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_17"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_17 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_17_r2),              
    .in_valid          (din_valid_4_17_r2),             
    .in_ready          (din_ready_4_17),             
    .out_data          (back_data_4_17),              
    .out_valid         (back_valid_4_17),             
    .out_ready         (back_ready_4_17),             
    .fill_level        (din_csr_readdata_4_17),
    .almost_full       (din_almost_full_4_17),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_18"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_18 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_18_r2),              
    .in_valid          (din_valid_4_18_r2),             
    .in_ready          (din_ready_4_18),             
    .out_data          (back_data_4_18),              
    .out_valid         (back_valid_4_18),             
    .out_ready         (back_ready_4_18),             
    .fill_level        (din_csr_readdata_4_18),
    .almost_full       (din_almost_full_4_18),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_19"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_19 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_19_r2),              
    .in_valid          (din_valid_4_19_r2),             
    .in_ready          (din_ready_4_19),             
    .out_data          (back_data_4_19),              
    .out_valid         (back_valid_4_19),             
    .out_ready         (back_ready_4_19),             
    .fill_level        (din_csr_readdata_4_19),
    .almost_full       (din_almost_full_4_19),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_20"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_20 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_20_r2),              
    .in_valid          (din_valid_4_20_r2),             
    .in_ready          (din_ready_4_20),             
    .out_data          (back_data_4_20),              
    .out_valid         (back_valid_4_20),             
    .out_ready         (back_ready_4_20),             
    .fill_level        (din_csr_readdata_4_20),
    .almost_full       (din_almost_full_4_20),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_21"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_21 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_21_r2),              
    .in_valid          (din_valid_4_21_r2),             
    .in_ready          (din_ready_4_21),             
    .out_data          (back_data_4_21),              
    .out_valid         (back_valid_4_21),             
    .out_ready         (back_ready_4_21),             
    .fill_level        (din_csr_readdata_4_21),
    .almost_full       (din_almost_full_4_21),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_22"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_22 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_22_r2),              
    .in_valid          (din_valid_4_22_r2),             
    .in_ready          (din_ready_4_22),             
    .out_data          (back_data_4_22),              
    .out_valid         (back_valid_4_22),             
    .out_ready         (back_ready_4_22),             
    .fill_level        (din_csr_readdata_4_22),
    .almost_full       (din_almost_full_4_22),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_23"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_23 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_23_r2),              
    .in_valid          (din_valid_4_23_r2),             
    .in_ready          (din_ready_4_23),             
    .out_data          (back_data_4_23),              
    .out_valid         (back_valid_4_23),             
    .out_ready         (back_ready_4_23),             
    .fill_level        (din_csr_readdata_4_23),
    .almost_full       (din_almost_full_4_23),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_24"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_24 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_24_r2),              
    .in_valid          (din_valid_4_24_r2),             
    .in_ready          (din_ready_4_24),             
    .out_data          (back_data_4_24),              
    .out_valid         (back_valid_4_24),             
    .out_ready         (back_ready_4_24),             
    .fill_level        (din_csr_readdata_4_24),
    .almost_full       (din_almost_full_4_24),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_25"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_25 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_25_r2),              
    .in_valid          (din_valid_4_25_r2),             
    .in_ready          (din_ready_4_25),             
    .out_data          (back_data_4_25),              
    .out_valid         (back_valid_4_25),             
    .out_ready         (back_ready_4_25),             
    .fill_level        (din_csr_readdata_4_25),
    .almost_full       (din_almost_full_4_25),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_26"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_26 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_26_r2),              
    .in_valid          (din_valid_4_26_r2),             
    .in_ready          (din_ready_4_26),             
    .out_data          (back_data_4_26),              
    .out_valid         (back_valid_4_26),             
    .out_ready         (back_ready_4_26),             
    .fill_level        (din_csr_readdata_4_26),
    .almost_full       (din_almost_full_4_26),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_27"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_27 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_27_r2),              
    .in_valid          (din_valid_4_27_r2),             
    .in_ready          (din_ready_4_27),             
    .out_data          (back_data_4_27),              
    .out_valid         (back_valid_4_27),             
    .out_ready         (back_ready_4_27),             
    .fill_level        (din_csr_readdata_4_27),
    .almost_full       (din_almost_full_4_27),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_28"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_28 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_28_r2),              
    .in_valid          (din_valid_4_28_r2),             
    .in_ready          (din_ready_4_28),             
    .out_data          (back_data_4_28),              
    .out_valid         (back_valid_4_28),             
    .out_ready         (back_ready_4_28),             
    .fill_level        (din_csr_readdata_4_28),
    .almost_full       (din_almost_full_4_28),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_29"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_29 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_29_r2),              
    .in_valid          (din_valid_4_29_r2),             
    .in_ready          (din_ready_4_29),             
    .out_data          (back_data_4_29),              
    .out_valid         (back_valid_4_29),             
    .out_ready         (back_ready_4_29),             
    .fill_level        (din_csr_readdata_4_29),
    .almost_full       (din_almost_full_4_29),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_30"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_30 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_30_r2),              
    .in_valid          (din_valid_4_30_r2),             
    .in_ready          (din_ready_4_30),             
    .out_data          (back_data_4_30),              
    .out_valid         (back_valid_4_30),             
    .out_ready         (back_ready_4_30),             
    .fill_level        (din_csr_readdata_4_30),
    .almost_full       (din_almost_full_4_30),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_4_31"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_4_31 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_4_31_r2),              
    .in_valid          (din_valid_4_31_r2),             
    .in_ready          (din_ready_4_31),             
    .out_data          (back_data_4_31),              
    .out_valid         (back_valid_4_31),             
    .out_ready         (back_ready_4_31),             
    .fill_level        (din_csr_readdata_4_31),
    .almost_full       (din_almost_full_4_31),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_0"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_0 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_0_r2),              
    .in_valid          (din_valid_5_0_r2),             
    .in_ready          (din_ready_5_0),             
    .out_data          (back_data_5_0),              
    .out_valid         (back_valid_5_0),             
    .out_ready         (back_ready_5_0),             
    .fill_level        (din_csr_readdata_5_0),
    .almost_full       (din_almost_full_5_0),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_1"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_1 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_1_r2),              
    .in_valid          (din_valid_5_1_r2),             
    .in_ready          (din_ready_5_1),             
    .out_data          (back_data_5_1),              
    .out_valid         (back_valid_5_1),             
    .out_ready         (back_ready_5_1),             
    .fill_level        (din_csr_readdata_5_1),
    .almost_full       (din_almost_full_5_1),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_2"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_2 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_2_r2),              
    .in_valid          (din_valid_5_2_r2),             
    .in_ready          (din_ready_5_2),             
    .out_data          (back_data_5_2),              
    .out_valid         (back_valid_5_2),             
    .out_ready         (back_ready_5_2),             
    .fill_level        (din_csr_readdata_5_2),
    .almost_full       (din_almost_full_5_2),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_3"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_3 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_3_r2),              
    .in_valid          (din_valid_5_3_r2),             
    .in_ready          (din_ready_5_3),             
    .out_data          (back_data_5_3),              
    .out_valid         (back_valid_5_3),             
    .out_ready         (back_ready_5_3),             
    .fill_level        (din_csr_readdata_5_3),
    .almost_full       (din_almost_full_5_3),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_4"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_4 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_4_r2),              
    .in_valid          (din_valid_5_4_r2),             
    .in_ready          (din_ready_5_4),             
    .out_data          (back_data_5_4),              
    .out_valid         (back_valid_5_4),             
    .out_ready         (back_ready_5_4),             
    .fill_level        (din_csr_readdata_5_4),
    .almost_full       (din_almost_full_5_4),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_5"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_5 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_5_r2),              
    .in_valid          (din_valid_5_5_r2),             
    .in_ready          (din_ready_5_5),             
    .out_data          (back_data_5_5),              
    .out_valid         (back_valid_5_5),             
    .out_ready         (back_ready_5_5),             
    .fill_level        (din_csr_readdata_5_5),
    .almost_full       (din_almost_full_5_5),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_6"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_6 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_6_r2),              
    .in_valid          (din_valid_5_6_r2),             
    .in_ready          (din_ready_5_6),             
    .out_data          (back_data_5_6),              
    .out_valid         (back_valid_5_6),             
    .out_ready         (back_ready_5_6),             
    .fill_level        (din_csr_readdata_5_6),
    .almost_full       (din_almost_full_5_6),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_7"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_7 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_7_r2),              
    .in_valid          (din_valid_5_7_r2),             
    .in_ready          (din_ready_5_7),             
    .out_data          (back_data_5_7),              
    .out_valid         (back_valid_5_7),             
    .out_ready         (back_ready_5_7),             
    .fill_level        (din_csr_readdata_5_7),
    .almost_full       (din_almost_full_5_7),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_8"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_8 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_8_r2),              
    .in_valid          (din_valid_5_8_r2),             
    .in_ready          (din_ready_5_8),             
    .out_data          (back_data_5_8),              
    .out_valid         (back_valid_5_8),             
    .out_ready         (back_ready_5_8),             
    .fill_level        (din_csr_readdata_5_8),
    .almost_full       (din_almost_full_5_8),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_9"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_9 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_9_r2),              
    .in_valid          (din_valid_5_9_r2),             
    .in_ready          (din_ready_5_9),             
    .out_data          (back_data_5_9),              
    .out_valid         (back_valid_5_9),             
    .out_ready         (back_ready_5_9),             
    .fill_level        (din_csr_readdata_5_9),
    .almost_full       (din_almost_full_5_9),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_10"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_10 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_10_r2),              
    .in_valid          (din_valid_5_10_r2),             
    .in_ready          (din_ready_5_10),             
    .out_data          (back_data_5_10),              
    .out_valid         (back_valid_5_10),             
    .out_ready         (back_ready_5_10),             
    .fill_level        (din_csr_readdata_5_10),
    .almost_full       (din_almost_full_5_10),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_11"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_11 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_11_r2),              
    .in_valid          (din_valid_5_11_r2),             
    .in_ready          (din_ready_5_11),             
    .out_data          (back_data_5_11),              
    .out_valid         (back_valid_5_11),             
    .out_ready         (back_ready_5_11),             
    .fill_level        (din_csr_readdata_5_11),
    .almost_full       (din_almost_full_5_11),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_12"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_12 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_12_r2),              
    .in_valid          (din_valid_5_12_r2),             
    .in_ready          (din_ready_5_12),             
    .out_data          (back_data_5_12),              
    .out_valid         (back_valid_5_12),             
    .out_ready         (back_ready_5_12),             
    .fill_level        (din_csr_readdata_5_12),
    .almost_full       (din_almost_full_5_12),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_13"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_13 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_13_r2),              
    .in_valid          (din_valid_5_13_r2),             
    .in_ready          (din_ready_5_13),             
    .out_data          (back_data_5_13),              
    .out_valid         (back_valid_5_13),             
    .out_ready         (back_ready_5_13),             
    .fill_level        (din_csr_readdata_5_13),
    .almost_full       (din_almost_full_5_13),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_14"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_14 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_14_r2),              
    .in_valid          (din_valid_5_14_r2),             
    .in_ready          (din_ready_5_14),             
    .out_data          (back_data_5_14),              
    .out_valid         (back_valid_5_14),             
    .out_ready         (back_ready_5_14),             
    .fill_level        (din_csr_readdata_5_14),
    .almost_full       (din_almost_full_5_14),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_15"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_15 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_15_r2),              
    .in_valid          (din_valid_5_15_r2),             
    .in_ready          (din_ready_5_15),             
    .out_data          (back_data_5_15),              
    .out_valid         (back_valid_5_15),             
    .out_ready         (back_ready_5_15),             
    .fill_level        (din_csr_readdata_5_15),
    .almost_full       (din_almost_full_5_15),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_16"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_16 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_16_r2),              
    .in_valid          (din_valid_5_16_r2),             
    .in_ready          (din_ready_5_16),             
    .out_data          (back_data_5_16),              
    .out_valid         (back_valid_5_16),             
    .out_ready         (back_ready_5_16),             
    .fill_level        (din_csr_readdata_5_16),
    .almost_full       (din_almost_full_5_16),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_17"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_17 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_17_r2),              
    .in_valid          (din_valid_5_17_r2),             
    .in_ready          (din_ready_5_17),             
    .out_data          (back_data_5_17),              
    .out_valid         (back_valid_5_17),             
    .out_ready         (back_ready_5_17),             
    .fill_level        (din_csr_readdata_5_17),
    .almost_full       (din_almost_full_5_17),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_18"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_18 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_18_r2),              
    .in_valid          (din_valid_5_18_r2),             
    .in_ready          (din_ready_5_18),             
    .out_data          (back_data_5_18),              
    .out_valid         (back_valid_5_18),             
    .out_ready         (back_ready_5_18),             
    .fill_level        (din_csr_readdata_5_18),
    .almost_full       (din_almost_full_5_18),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_19"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_19 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_19_r2),              
    .in_valid          (din_valid_5_19_r2),             
    .in_ready          (din_ready_5_19),             
    .out_data          (back_data_5_19),              
    .out_valid         (back_valid_5_19),             
    .out_ready         (back_ready_5_19),             
    .fill_level        (din_csr_readdata_5_19),
    .almost_full       (din_almost_full_5_19),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_20"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_20 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_20_r2),              
    .in_valid          (din_valid_5_20_r2),             
    .in_ready          (din_ready_5_20),             
    .out_data          (back_data_5_20),              
    .out_valid         (back_valid_5_20),             
    .out_ready         (back_ready_5_20),             
    .fill_level        (din_csr_readdata_5_20),
    .almost_full       (din_almost_full_5_20),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_21"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_21 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_21_r2),              
    .in_valid          (din_valid_5_21_r2),             
    .in_ready          (din_ready_5_21),             
    .out_data          (back_data_5_21),              
    .out_valid         (back_valid_5_21),             
    .out_ready         (back_ready_5_21),             
    .fill_level        (din_csr_readdata_5_21),
    .almost_full       (din_almost_full_5_21),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_22"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_22 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_22_r2),              
    .in_valid          (din_valid_5_22_r2),             
    .in_ready          (din_ready_5_22),             
    .out_data          (back_data_5_22),              
    .out_valid         (back_valid_5_22),             
    .out_ready         (back_ready_5_22),             
    .fill_level        (din_csr_readdata_5_22),
    .almost_full       (din_almost_full_5_22),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_23"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_23 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_23_r2),              
    .in_valid          (din_valid_5_23_r2),             
    .in_ready          (din_ready_5_23),             
    .out_data          (back_data_5_23),              
    .out_valid         (back_valid_5_23),             
    .out_ready         (back_ready_5_23),             
    .fill_level        (din_csr_readdata_5_23),
    .almost_full       (din_almost_full_5_23),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_24"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_24 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_24_r2),              
    .in_valid          (din_valid_5_24_r2),             
    .in_ready          (din_ready_5_24),             
    .out_data          (back_data_5_24),              
    .out_valid         (back_valid_5_24),             
    .out_ready         (back_ready_5_24),             
    .fill_level        (din_csr_readdata_5_24),
    .almost_full       (din_almost_full_5_24),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_25"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_25 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_25_r2),              
    .in_valid          (din_valid_5_25_r2),             
    .in_ready          (din_ready_5_25),             
    .out_data          (back_data_5_25),              
    .out_valid         (back_valid_5_25),             
    .out_ready         (back_ready_5_25),             
    .fill_level        (din_csr_readdata_5_25),
    .almost_full       (din_almost_full_5_25),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_26"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_26 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_26_r2),              
    .in_valid          (din_valid_5_26_r2),             
    .in_ready          (din_ready_5_26),             
    .out_data          (back_data_5_26),              
    .out_valid         (back_valid_5_26),             
    .out_ready         (back_ready_5_26),             
    .fill_level        (din_csr_readdata_5_26),
    .almost_full       (din_almost_full_5_26),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_27"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_27 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_27_r2),              
    .in_valid          (din_valid_5_27_r2),             
    .in_ready          (din_ready_5_27),             
    .out_data          (back_data_5_27),              
    .out_valid         (back_valid_5_27),             
    .out_ready         (back_ready_5_27),             
    .fill_level        (din_csr_readdata_5_27),
    .almost_full       (din_almost_full_5_27),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_28"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_28 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_28_r2),              
    .in_valid          (din_valid_5_28_r2),             
    .in_ready          (din_ready_5_28),             
    .out_data          (back_data_5_28),              
    .out_valid         (back_valid_5_28),             
    .out_ready         (back_ready_5_28),             
    .fill_level        (din_csr_readdata_5_28),
    .almost_full       (din_almost_full_5_28),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_29"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_29 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_29_r2),              
    .in_valid          (din_valid_5_29_r2),             
    .in_ready          (din_ready_5_29),             
    .out_data          (back_data_5_29),              
    .out_valid         (back_valid_5_29),             
    .out_ready         (back_ready_5_29),             
    .fill_level        (din_csr_readdata_5_29),
    .almost_full       (din_almost_full_5_29),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_30"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_30 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_30_r2),              
    .in_valid          (din_valid_5_30_r2),             
    .in_ready          (din_ready_5_30),             
    .out_data          (back_data_5_30),              
    .out_valid         (back_valid_5_30),             
    .out_ready         (back_ready_5_30),             
    .fill_level        (din_csr_readdata_5_30),
    .almost_full       (din_almost_full_5_30),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_5_31"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_5_31 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_5_31_r2),              
    .in_valid          (din_valid_5_31_r2),             
    .in_ready          (din_ready_5_31),             
    .out_data          (back_data_5_31),              
    .out_valid         (back_valid_5_31),             
    .out_ready         (back_ready_5_31),             
    .fill_level        (din_csr_readdata_5_31),
    .almost_full       (din_almost_full_5_31),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_0"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_0 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_0_r2),              
    .in_valid          (din_valid_6_0_r2),             
    .in_ready          (din_ready_6_0),             
    .out_data          (back_data_6_0),              
    .out_valid         (back_valid_6_0),             
    .out_ready         (back_ready_6_0),             
    .fill_level        (din_csr_readdata_6_0),
    .almost_full       (din_almost_full_6_0),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_1"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_1 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_1_r2),              
    .in_valid          (din_valid_6_1_r2),             
    .in_ready          (din_ready_6_1),             
    .out_data          (back_data_6_1),              
    .out_valid         (back_valid_6_1),             
    .out_ready         (back_ready_6_1),             
    .fill_level        (din_csr_readdata_6_1),
    .almost_full       (din_almost_full_6_1),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_2"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_2 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_2_r2),              
    .in_valid          (din_valid_6_2_r2),             
    .in_ready          (din_ready_6_2),             
    .out_data          (back_data_6_2),              
    .out_valid         (back_valid_6_2),             
    .out_ready         (back_ready_6_2),             
    .fill_level        (din_csr_readdata_6_2),
    .almost_full       (din_almost_full_6_2),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_3"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_3 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_3_r2),              
    .in_valid          (din_valid_6_3_r2),             
    .in_ready          (din_ready_6_3),             
    .out_data          (back_data_6_3),              
    .out_valid         (back_valid_6_3),             
    .out_ready         (back_ready_6_3),             
    .fill_level        (din_csr_readdata_6_3),
    .almost_full       (din_almost_full_6_3),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_4"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_4 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_4_r2),              
    .in_valid          (din_valid_6_4_r2),             
    .in_ready          (din_ready_6_4),             
    .out_data          (back_data_6_4),              
    .out_valid         (back_valid_6_4),             
    .out_ready         (back_ready_6_4),             
    .fill_level        (din_csr_readdata_6_4),
    .almost_full       (din_almost_full_6_4),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_5"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_5 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_5_r2),              
    .in_valid          (din_valid_6_5_r2),             
    .in_ready          (din_ready_6_5),             
    .out_data          (back_data_6_5),              
    .out_valid         (back_valid_6_5),             
    .out_ready         (back_ready_6_5),             
    .fill_level        (din_csr_readdata_6_5),
    .almost_full       (din_almost_full_6_5),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_6"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_6 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_6_r2),              
    .in_valid          (din_valid_6_6_r2),             
    .in_ready          (din_ready_6_6),             
    .out_data          (back_data_6_6),              
    .out_valid         (back_valid_6_6),             
    .out_ready         (back_ready_6_6),             
    .fill_level        (din_csr_readdata_6_6),
    .almost_full       (din_almost_full_6_6),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_7"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_7 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_7_r2),              
    .in_valid          (din_valid_6_7_r2),             
    .in_ready          (din_ready_6_7),             
    .out_data          (back_data_6_7),              
    .out_valid         (back_valid_6_7),             
    .out_ready         (back_ready_6_7),             
    .fill_level        (din_csr_readdata_6_7),
    .almost_full       (din_almost_full_6_7),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_8"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_8 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_8_r2),              
    .in_valid          (din_valid_6_8_r2),             
    .in_ready          (din_ready_6_8),             
    .out_data          (back_data_6_8),              
    .out_valid         (back_valid_6_8),             
    .out_ready         (back_ready_6_8),             
    .fill_level        (din_csr_readdata_6_8),
    .almost_full       (din_almost_full_6_8),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_9"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_9 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_9_r2),              
    .in_valid          (din_valid_6_9_r2),             
    .in_ready          (din_ready_6_9),             
    .out_data          (back_data_6_9),              
    .out_valid         (back_valid_6_9),             
    .out_ready         (back_ready_6_9),             
    .fill_level        (din_csr_readdata_6_9),
    .almost_full       (din_almost_full_6_9),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_10"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_10 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_10_r2),              
    .in_valid          (din_valid_6_10_r2),             
    .in_ready          (din_ready_6_10),             
    .out_data          (back_data_6_10),              
    .out_valid         (back_valid_6_10),             
    .out_ready         (back_ready_6_10),             
    .fill_level        (din_csr_readdata_6_10),
    .almost_full       (din_almost_full_6_10),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_11"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_11 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_11_r2),              
    .in_valid          (din_valid_6_11_r2),             
    .in_ready          (din_ready_6_11),             
    .out_data          (back_data_6_11),              
    .out_valid         (back_valid_6_11),             
    .out_ready         (back_ready_6_11),             
    .fill_level        (din_csr_readdata_6_11),
    .almost_full       (din_almost_full_6_11),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_12"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_12 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_12_r2),              
    .in_valid          (din_valid_6_12_r2),             
    .in_ready          (din_ready_6_12),             
    .out_data          (back_data_6_12),              
    .out_valid         (back_valid_6_12),             
    .out_ready         (back_ready_6_12),             
    .fill_level        (din_csr_readdata_6_12),
    .almost_full       (din_almost_full_6_12),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_13"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_13 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_13_r2),              
    .in_valid          (din_valid_6_13_r2),             
    .in_ready          (din_ready_6_13),             
    .out_data          (back_data_6_13),              
    .out_valid         (back_valid_6_13),             
    .out_ready         (back_ready_6_13),             
    .fill_level        (din_csr_readdata_6_13),
    .almost_full       (din_almost_full_6_13),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_14"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_14 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_14_r2),              
    .in_valid          (din_valid_6_14_r2),             
    .in_ready          (din_ready_6_14),             
    .out_data          (back_data_6_14),              
    .out_valid         (back_valid_6_14),             
    .out_ready         (back_ready_6_14),             
    .fill_level        (din_csr_readdata_6_14),
    .almost_full       (din_almost_full_6_14),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_15"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_15 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_15_r2),              
    .in_valid          (din_valid_6_15_r2),             
    .in_ready          (din_ready_6_15),             
    .out_data          (back_data_6_15),              
    .out_valid         (back_valid_6_15),             
    .out_ready         (back_ready_6_15),             
    .fill_level        (din_csr_readdata_6_15),
    .almost_full       (din_almost_full_6_15),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_16"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_16 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_16_r2),              
    .in_valid          (din_valid_6_16_r2),             
    .in_ready          (din_ready_6_16),             
    .out_data          (back_data_6_16),              
    .out_valid         (back_valid_6_16),             
    .out_ready         (back_ready_6_16),             
    .fill_level        (din_csr_readdata_6_16),
    .almost_full       (din_almost_full_6_16),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_17"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_17 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_17_r2),              
    .in_valid          (din_valid_6_17_r2),             
    .in_ready          (din_ready_6_17),             
    .out_data          (back_data_6_17),              
    .out_valid         (back_valid_6_17),             
    .out_ready         (back_ready_6_17),             
    .fill_level        (din_csr_readdata_6_17),
    .almost_full       (din_almost_full_6_17),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_18"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_18 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_18_r2),              
    .in_valid          (din_valid_6_18_r2),             
    .in_ready          (din_ready_6_18),             
    .out_data          (back_data_6_18),              
    .out_valid         (back_valid_6_18),             
    .out_ready         (back_ready_6_18),             
    .fill_level        (din_csr_readdata_6_18),
    .almost_full       (din_almost_full_6_18),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_19"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_19 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_19_r2),              
    .in_valid          (din_valid_6_19_r2),             
    .in_ready          (din_ready_6_19),             
    .out_data          (back_data_6_19),              
    .out_valid         (back_valid_6_19),             
    .out_ready         (back_ready_6_19),             
    .fill_level        (din_csr_readdata_6_19),
    .almost_full       (din_almost_full_6_19),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_20"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_20 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_20_r2),              
    .in_valid          (din_valid_6_20_r2),             
    .in_ready          (din_ready_6_20),             
    .out_data          (back_data_6_20),              
    .out_valid         (back_valid_6_20),             
    .out_ready         (back_ready_6_20),             
    .fill_level        (din_csr_readdata_6_20),
    .almost_full       (din_almost_full_6_20),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_21"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_21 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_21_r2),              
    .in_valid          (din_valid_6_21_r2),             
    .in_ready          (din_ready_6_21),             
    .out_data          (back_data_6_21),              
    .out_valid         (back_valid_6_21),             
    .out_ready         (back_ready_6_21),             
    .fill_level        (din_csr_readdata_6_21),
    .almost_full       (din_almost_full_6_21),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_22"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_22 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_22_r2),              
    .in_valid          (din_valid_6_22_r2),             
    .in_ready          (din_ready_6_22),             
    .out_data          (back_data_6_22),              
    .out_valid         (back_valid_6_22),             
    .out_ready         (back_ready_6_22),             
    .fill_level        (din_csr_readdata_6_22),
    .almost_full       (din_almost_full_6_22),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_23"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_23 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_23_r2),              
    .in_valid          (din_valid_6_23_r2),             
    .in_ready          (din_ready_6_23),             
    .out_data          (back_data_6_23),              
    .out_valid         (back_valid_6_23),             
    .out_ready         (back_ready_6_23),             
    .fill_level        (din_csr_readdata_6_23),
    .almost_full       (din_almost_full_6_23),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_24"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_24 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_24_r2),              
    .in_valid          (din_valid_6_24_r2),             
    .in_ready          (din_ready_6_24),             
    .out_data          (back_data_6_24),              
    .out_valid         (back_valid_6_24),             
    .out_ready         (back_ready_6_24),             
    .fill_level        (din_csr_readdata_6_24),
    .almost_full       (din_almost_full_6_24),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_25"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_25 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_25_r2),              
    .in_valid          (din_valid_6_25_r2),             
    .in_ready          (din_ready_6_25),             
    .out_data          (back_data_6_25),              
    .out_valid         (back_valid_6_25),             
    .out_ready         (back_ready_6_25),             
    .fill_level        (din_csr_readdata_6_25),
    .almost_full       (din_almost_full_6_25),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_26"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_26 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_26_r2),              
    .in_valid          (din_valid_6_26_r2),             
    .in_ready          (din_ready_6_26),             
    .out_data          (back_data_6_26),              
    .out_valid         (back_valid_6_26),             
    .out_ready         (back_ready_6_26),             
    .fill_level        (din_csr_readdata_6_26),
    .almost_full       (din_almost_full_6_26),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_27"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_27 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_27_r2),              
    .in_valid          (din_valid_6_27_r2),             
    .in_ready          (din_ready_6_27),             
    .out_data          (back_data_6_27),              
    .out_valid         (back_valid_6_27),             
    .out_ready         (back_ready_6_27),             
    .fill_level        (din_csr_readdata_6_27),
    .almost_full       (din_almost_full_6_27),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_28"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_28 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_28_r2),              
    .in_valid          (din_valid_6_28_r2),             
    .in_ready          (din_ready_6_28),             
    .out_data          (back_data_6_28),              
    .out_valid         (back_valid_6_28),             
    .out_ready         (back_ready_6_28),             
    .fill_level        (din_csr_readdata_6_28),
    .almost_full       (din_almost_full_6_28),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_29"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_29 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_29_r2),              
    .in_valid          (din_valid_6_29_r2),             
    .in_ready          (din_ready_6_29),             
    .out_data          (back_data_6_29),              
    .out_valid         (back_valid_6_29),             
    .out_ready         (back_ready_6_29),             
    .fill_level        (din_csr_readdata_6_29),
    .almost_full       (din_almost_full_6_29),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_30"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_30 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_30_r2),              
    .in_valid          (din_valid_6_30_r2),             
    .in_ready          (din_ready_6_30),             
    .out_data          (back_data_6_30),              
    .out_valid         (back_valid_6_30),             
    .out_ready         (back_ready_6_30),             
    .fill_level        (din_csr_readdata_6_30),
    .almost_full       (din_almost_full_6_30),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_6_31"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_6_31 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_6_31_r2),              
    .in_valid          (din_valid_6_31_r2),             
    .in_ready          (din_ready_6_31),             
    .out_data          (back_data_6_31),              
    .out_valid         (back_valid_6_31),             
    .out_ready         (back_ready_6_31),             
    .fill_level        (din_csr_readdata_6_31),
    .almost_full       (din_almost_full_6_31),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_0"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_0 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_0_r2),              
    .in_valid          (din_valid_7_0_r2),             
    .in_ready          (din_ready_7_0),             
    .out_data          (back_data_7_0),              
    .out_valid         (back_valid_7_0),             
    .out_ready         (back_ready_7_0),             
    .fill_level        (din_csr_readdata_7_0),
    .almost_full       (din_almost_full_7_0),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_1"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_1 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_1_r2),              
    .in_valid          (din_valid_7_1_r2),             
    .in_ready          (din_ready_7_1),             
    .out_data          (back_data_7_1),              
    .out_valid         (back_valid_7_1),             
    .out_ready         (back_ready_7_1),             
    .fill_level        (din_csr_readdata_7_1),
    .almost_full       (din_almost_full_7_1),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_2"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_2 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_2_r2),              
    .in_valid          (din_valid_7_2_r2),             
    .in_ready          (din_ready_7_2),             
    .out_data          (back_data_7_2),              
    .out_valid         (back_valid_7_2),             
    .out_ready         (back_ready_7_2),             
    .fill_level        (din_csr_readdata_7_2),
    .almost_full       (din_almost_full_7_2),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_3"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_3 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_3_r2),              
    .in_valid          (din_valid_7_3_r2),             
    .in_ready          (din_ready_7_3),             
    .out_data          (back_data_7_3),              
    .out_valid         (back_valid_7_3),             
    .out_ready         (back_ready_7_3),             
    .fill_level        (din_csr_readdata_7_3),
    .almost_full       (din_almost_full_7_3),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_4"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_4 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_4_r2),              
    .in_valid          (din_valid_7_4_r2),             
    .in_ready          (din_ready_7_4),             
    .out_data          (back_data_7_4),              
    .out_valid         (back_valid_7_4),             
    .out_ready         (back_ready_7_4),             
    .fill_level        (din_csr_readdata_7_4),
    .almost_full       (din_almost_full_7_4),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_5"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_5 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_5_r2),              
    .in_valid          (din_valid_7_5_r2),             
    .in_ready          (din_ready_7_5),             
    .out_data          (back_data_7_5),              
    .out_valid         (back_valid_7_5),             
    .out_ready         (back_ready_7_5),             
    .fill_level        (din_csr_readdata_7_5),
    .almost_full       (din_almost_full_7_5),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_6"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_6 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_6_r2),              
    .in_valid          (din_valid_7_6_r2),             
    .in_ready          (din_ready_7_6),             
    .out_data          (back_data_7_6),              
    .out_valid         (back_valid_7_6),             
    .out_ready         (back_ready_7_6),             
    .fill_level        (din_csr_readdata_7_6),
    .almost_full       (din_almost_full_7_6),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_7"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_7 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_7_r2),              
    .in_valid          (din_valid_7_7_r2),             
    .in_ready          (din_ready_7_7),             
    .out_data          (back_data_7_7),              
    .out_valid         (back_valid_7_7),             
    .out_ready         (back_ready_7_7),             
    .fill_level        (din_csr_readdata_7_7),
    .almost_full       (din_almost_full_7_7),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_8"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_8 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_8_r2),              
    .in_valid          (din_valid_7_8_r2),             
    .in_ready          (din_ready_7_8),             
    .out_data          (back_data_7_8),              
    .out_valid         (back_valid_7_8),             
    .out_ready         (back_ready_7_8),             
    .fill_level        (din_csr_readdata_7_8),
    .almost_full       (din_almost_full_7_8),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_9"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_9 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_9_r2),              
    .in_valid          (din_valid_7_9_r2),             
    .in_ready          (din_ready_7_9),             
    .out_data          (back_data_7_9),              
    .out_valid         (back_valid_7_9),             
    .out_ready         (back_ready_7_9),             
    .fill_level        (din_csr_readdata_7_9),
    .almost_full       (din_almost_full_7_9),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_10"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_10 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_10_r2),              
    .in_valid          (din_valid_7_10_r2),             
    .in_ready          (din_ready_7_10),             
    .out_data          (back_data_7_10),              
    .out_valid         (back_valid_7_10),             
    .out_ready         (back_ready_7_10),             
    .fill_level        (din_csr_readdata_7_10),
    .almost_full       (din_almost_full_7_10),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_11"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_11 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_11_r2),              
    .in_valid          (din_valid_7_11_r2),             
    .in_ready          (din_ready_7_11),             
    .out_data          (back_data_7_11),              
    .out_valid         (back_valid_7_11),             
    .out_ready         (back_ready_7_11),             
    .fill_level        (din_csr_readdata_7_11),
    .almost_full       (din_almost_full_7_11),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_12"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_12 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_12_r2),              
    .in_valid          (din_valid_7_12_r2),             
    .in_ready          (din_ready_7_12),             
    .out_data          (back_data_7_12),              
    .out_valid         (back_valid_7_12),             
    .out_ready         (back_ready_7_12),             
    .fill_level        (din_csr_readdata_7_12),
    .almost_full       (din_almost_full_7_12),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_13"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_13 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_13_r2),              
    .in_valid          (din_valid_7_13_r2),             
    .in_ready          (din_ready_7_13),             
    .out_data          (back_data_7_13),              
    .out_valid         (back_valid_7_13),             
    .out_ready         (back_ready_7_13),             
    .fill_level        (din_csr_readdata_7_13),
    .almost_full       (din_almost_full_7_13),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_14"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_14 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_14_r2),              
    .in_valid          (din_valid_7_14_r2),             
    .in_ready          (din_ready_7_14),             
    .out_data          (back_data_7_14),              
    .out_valid         (back_valid_7_14),             
    .out_ready         (back_ready_7_14),             
    .fill_level        (din_csr_readdata_7_14),
    .almost_full       (din_almost_full_7_14),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_15"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_15 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_15_r2),              
    .in_valid          (din_valid_7_15_r2),             
    .in_ready          (din_ready_7_15),             
    .out_data          (back_data_7_15),              
    .out_valid         (back_valid_7_15),             
    .out_ready         (back_ready_7_15),             
    .fill_level        (din_csr_readdata_7_15),
    .almost_full       (din_almost_full_7_15),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_16"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_16 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_16_r2),              
    .in_valid          (din_valid_7_16_r2),             
    .in_ready          (din_ready_7_16),             
    .out_data          (back_data_7_16),              
    .out_valid         (back_valid_7_16),             
    .out_ready         (back_ready_7_16),             
    .fill_level        (din_csr_readdata_7_16),
    .almost_full       (din_almost_full_7_16),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_17"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_17 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_17_r2),              
    .in_valid          (din_valid_7_17_r2),             
    .in_ready          (din_ready_7_17),             
    .out_data          (back_data_7_17),              
    .out_valid         (back_valid_7_17),             
    .out_ready         (back_ready_7_17),             
    .fill_level        (din_csr_readdata_7_17),
    .almost_full       (din_almost_full_7_17),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_18"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_18 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_18_r2),              
    .in_valid          (din_valid_7_18_r2),             
    .in_ready          (din_ready_7_18),             
    .out_data          (back_data_7_18),              
    .out_valid         (back_valid_7_18),             
    .out_ready         (back_ready_7_18),             
    .fill_level        (din_csr_readdata_7_18),
    .almost_full       (din_almost_full_7_18),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_19"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_19 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_19_r2),              
    .in_valid          (din_valid_7_19_r2),             
    .in_ready          (din_ready_7_19),             
    .out_data          (back_data_7_19),              
    .out_valid         (back_valid_7_19),             
    .out_ready         (back_ready_7_19),             
    .fill_level        (din_csr_readdata_7_19),
    .almost_full       (din_almost_full_7_19),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_20"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_20 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_20_r2),              
    .in_valid          (din_valid_7_20_r2),             
    .in_ready          (din_ready_7_20),             
    .out_data          (back_data_7_20),              
    .out_valid         (back_valid_7_20),             
    .out_ready         (back_ready_7_20),             
    .fill_level        (din_csr_readdata_7_20),
    .almost_full       (din_almost_full_7_20),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_21"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_21 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_21_r2),              
    .in_valid          (din_valid_7_21_r2),             
    .in_ready          (din_ready_7_21),             
    .out_data          (back_data_7_21),              
    .out_valid         (back_valid_7_21),             
    .out_ready         (back_ready_7_21),             
    .fill_level        (din_csr_readdata_7_21),
    .almost_full       (din_almost_full_7_21),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_22"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_22 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_22_r2),              
    .in_valid          (din_valid_7_22_r2),             
    .in_ready          (din_ready_7_22),             
    .out_data          (back_data_7_22),              
    .out_valid         (back_valid_7_22),             
    .out_ready         (back_ready_7_22),             
    .fill_level        (din_csr_readdata_7_22),
    .almost_full       (din_almost_full_7_22),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_23"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_23 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_23_r2),              
    .in_valid          (din_valid_7_23_r2),             
    .in_ready          (din_ready_7_23),             
    .out_data          (back_data_7_23),              
    .out_valid         (back_valid_7_23),             
    .out_ready         (back_ready_7_23),             
    .fill_level        (din_csr_readdata_7_23),
    .almost_full       (din_almost_full_7_23),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_24"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_24 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_24_r2),              
    .in_valid          (din_valid_7_24_r2),             
    .in_ready          (din_ready_7_24),             
    .out_data          (back_data_7_24),              
    .out_valid         (back_valid_7_24),             
    .out_ready         (back_ready_7_24),             
    .fill_level        (din_csr_readdata_7_24),
    .almost_full       (din_almost_full_7_24),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_25"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_25 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_25_r2),              
    .in_valid          (din_valid_7_25_r2),             
    .in_ready          (din_ready_7_25),             
    .out_data          (back_data_7_25),              
    .out_valid         (back_valid_7_25),             
    .out_ready         (back_ready_7_25),             
    .fill_level        (din_csr_readdata_7_25),
    .almost_full       (din_almost_full_7_25),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_26"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_26 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_26_r2),              
    .in_valid          (din_valid_7_26_r2),             
    .in_ready          (din_ready_7_26),             
    .out_data          (back_data_7_26),              
    .out_valid         (back_valid_7_26),             
    .out_ready         (back_ready_7_26),             
    .fill_level        (din_csr_readdata_7_26),
    .almost_full       (din_almost_full_7_26),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_27"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_27 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_27_r2),              
    .in_valid          (din_valid_7_27_r2),             
    .in_ready          (din_ready_7_27),             
    .out_data          (back_data_7_27),              
    .out_valid         (back_valid_7_27),             
    .out_ready         (back_ready_7_27),             
    .fill_level        (din_csr_readdata_7_27),
    .almost_full       (din_almost_full_7_27),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_28"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_28 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_28_r2),              
    .in_valid          (din_valid_7_28_r2),             
    .in_ready          (din_ready_7_28),             
    .out_data          (back_data_7_28),              
    .out_valid         (back_valid_7_28),             
    .out_ready         (back_ready_7_28),             
    .fill_level        (din_csr_readdata_7_28),
    .almost_full       (din_almost_full_7_28),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_29"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_29 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_29_r2),              
    .in_valid          (din_valid_7_29_r2),             
    .in_ready          (din_ready_7_29),             
    .out_data          (back_data_7_29),              
    .out_valid         (back_valid_7_29),             
    .out_ready         (back_ready_7_29),             
    .fill_level        (din_csr_readdata_7_29),
    .almost_full       (din_almost_full_7_29),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_30"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_30 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_30_r2),              
    .in_valid          (din_valid_7_30_r2),             
    .in_ready          (din_ready_7_30),             
    .out_data          (back_data_7_30),              
    .out_valid         (back_valid_7_30),             
    .out_ready         (back_ready_7_30),             
    .fill_level        (din_csr_readdata_7_30),
    .almost_full       (din_almost_full_7_30),
    .overflow          ()
);
unified_fifo  #(
    .FIFO_NAME        ("[fast_pattern] dc_FIFO_7_31"),
    .MEM_TYPE         ("MLAB"),
    .DUAL_CLOCK       (1),
    .USE_ALMOST_FULL  (1),
    .FULL_LEVEL       (40),
    .SYMBOLS_PER_BEAT (1),
    .BITS_PER_SYMBOL  (RULE_S_WIDTH),
    .FIFO_DEPTH       (128)
) l1_dc_fifo_mlab_7_31 (
    .in_clk            (front_clk),
    .in_reset          (front_rst),
    .out_clk           (back_clk),
    .out_reset         (back_rst),
    .in_data           (din_7_31_r2),              
    .in_valid          (din_valid_7_31_r2),             
    .in_ready          (din_ready_7_31),             
    .out_data          (back_data_7_31),              
    .out_valid         (back_valid_7_31),             
    .out_ready         (back_ready_7_31),             
    .fill_level        (din_csr_readdata_7_31),
    .almost_full       (din_almost_full_7_31),
    .overflow          ()
);

`endif

`ifdef DEBUG
stats_cnt_rule #(.DEBUG(1))
out_rule_inst(
    .Clk        (back_clk),
    .Rst_n      (!back_rst),
    .valid      (out_usr_valid),
    .ready      (out_usr_ready),
    .data       (out_usr_data),
    .eop        (out_usr_eop),
    .sop        (out_usr_sop),
    .stats_rule ()
);
`endif
	
endmodule
`include "./src/struct_s.sv"
module cal_fp(
    input clk,
    input rst,
    output logic [FP_WIDTH-1:0] fp_data,
    output logic                fp_valid,
    input [NF_WIDTH-1:0] din_0_0,
    input din_valid_0_0,
    input [NF_WIDTH-1:0] din_0_1,
    input din_valid_0_1,
    input [NF_WIDTH-1:0] din_0_2,
    input din_valid_0_2,
    input [NF_WIDTH-1:0] din_0_3,
    input din_valid_0_3,
    input [NF_WIDTH-1:0] din_0_4,
    input din_valid_0_4,
    input [NF_WIDTH-1:0] din_0_5,
    input din_valid_0_5,
    input [NF_WIDTH-1:0] din_0_6,
    input din_valid_0_6,
    input [NF_WIDTH-1:0] din_0_7,
    input din_valid_0_7,
    input [NF_WIDTH-1:0] din_0_8,
    input din_valid_0_8,
    input [NF_WIDTH-1:0] din_0_9,
    input din_valid_0_9,
    input [NF_WIDTH-1:0] din_0_10,
    input din_valid_0_10,
    input [NF_WIDTH-1:0] din_0_11,
    input din_valid_0_11,
    input [NF_WIDTH-1:0] din_0_12,
    input din_valid_0_12,
    input [NF_WIDTH-1:0] din_0_13,
    input din_valid_0_13,
    input [NF_WIDTH-1:0] din_0_14,
    input din_valid_0_14,
    input [NF_WIDTH-1:0] din_0_15,
    input din_valid_0_15,
    input [NF_WIDTH-1:0] din_1_0,
    input din_valid_1_0,
    input [NF_WIDTH-1:0] din_1_1,
    input din_valid_1_1,
    input [NF_WIDTH-1:0] din_1_2,
    input din_valid_1_2,
    input [NF_WIDTH-1:0] din_1_3,
    input din_valid_1_3,
    input [NF_WIDTH-1:0] din_1_4,
    input din_valid_1_4,
    input [NF_WIDTH-1:0] din_1_5,
    input din_valid_1_5,
    input [NF_WIDTH-1:0] din_1_6,
    input din_valid_1_6,
    input [NF_WIDTH-1:0] din_1_7,
    input din_valid_1_7,
    input [NF_WIDTH-1:0] din_1_8,
    input din_valid_1_8,
    input [NF_WIDTH-1:0] din_1_9,
    input din_valid_1_9,
    input [NF_WIDTH-1:0] din_1_10,
    input din_valid_1_10,
    input [NF_WIDTH-1:0] din_1_11,
    input din_valid_1_11,
    input [NF_WIDTH-1:0] din_1_12,
    input din_valid_1_12,
    input [NF_WIDTH-1:0] din_1_13,
    input din_valid_1_13,
    input [NF_WIDTH-1:0] din_1_14,
    input din_valid_1_14,
    input [NF_WIDTH-1:0] din_1_15,
    input din_valid_1_15,
    input [NF_WIDTH-1:0] din_2_0,
    input din_valid_2_0,
    input [NF_WIDTH-1:0] din_2_1,
    input din_valid_2_1,
    input [NF_WIDTH-1:0] din_2_2,
    input din_valid_2_2,
    input [NF_WIDTH-1:0] din_2_3,
    input din_valid_2_3,
    input [NF_WIDTH-1:0] din_2_4,
    input din_valid_2_4,
    input [NF_WIDTH-1:0] din_2_5,
    input din_valid_2_5,
    input [NF_WIDTH-1:0] din_2_6,
    input din_valid_2_6,
    input [NF_WIDTH-1:0] din_2_7,
    input din_valid_2_7,
    input [NF_WIDTH-1:0] din_2_8,
    input din_valid_2_8,
    input [NF_WIDTH-1:0] din_2_9,
    input din_valid_2_9,
    input [NF_WIDTH-1:0] din_2_10,
    input din_valid_2_10,
    input [NF_WIDTH-1:0] din_2_11,
    input din_valid_2_11,
    input [NF_WIDTH-1:0] din_2_12,
    input din_valid_2_12,
    input [NF_WIDTH-1:0] din_2_13,
    input din_valid_2_13,
    input [NF_WIDTH-1:0] din_2_14,
    input din_valid_2_14,
    input [NF_WIDTH-1:0] din_2_15,
    input din_valid_2_15,
    input [NF_WIDTH-1:0] din_3_0,
    input din_valid_3_0,
    input [NF_WIDTH-1:0] din_3_1,
    input din_valid_3_1,
    input [NF_WIDTH-1:0] din_3_2,
    input din_valid_3_2,
    input [NF_WIDTH-1:0] din_3_3,
    input din_valid_3_3,
    input [NF_WIDTH-1:0] din_3_4,
    input din_valid_3_4,
    input [NF_WIDTH-1:0] din_3_5,
    input din_valid_3_5,
    input [NF_WIDTH-1:0] din_3_6,
    input din_valid_3_6,
    input [NF_WIDTH-1:0] din_3_7,
    input din_valid_3_7,
    input [NF_WIDTH-1:0] din_3_8,
    input din_valid_3_8,
    input [NF_WIDTH-1:0] din_3_9,
    input din_valid_3_9,
    input [NF_WIDTH-1:0] din_3_10,
    input din_valid_3_10,
    input [NF_WIDTH-1:0] din_3_11,
    input din_valid_3_11,
    input [NF_WIDTH-1:0] din_3_12,
    input din_valid_3_12,
    input [NF_WIDTH-1:0] din_3_13,
    input din_valid_3_13,
    input [NF_WIDTH-1:0] din_3_14,
    input din_valid_3_14,
    input [NF_WIDTH-1:0] din_3_15,
    input din_valid_3_15,
    input [NF_WIDTH-1:0] din_4_0,
    input din_valid_4_0,
    input [NF_WIDTH-1:0] din_4_1,
    input din_valid_4_1,
    input [NF_WIDTH-1:0] din_4_2,
    input din_valid_4_2,
    input [NF_WIDTH-1:0] din_4_3,
    input din_valid_4_3,
    input [NF_WIDTH-1:0] din_4_4,
    input din_valid_4_4,
    input [NF_WIDTH-1:0] din_4_5,
    input din_valid_4_5,
    input [NF_WIDTH-1:0] din_4_6,
    input din_valid_4_6,
    input [NF_WIDTH-1:0] din_4_7,
    input din_valid_4_7,
    input [NF_WIDTH-1:0] din_4_8,
    input din_valid_4_8,
    input [NF_WIDTH-1:0] din_4_9,
    input din_valid_4_9,
    input [NF_WIDTH-1:0] din_4_10,
    input din_valid_4_10,
    input [NF_WIDTH-1:0] din_4_11,
    input din_valid_4_11,
    input [NF_WIDTH-1:0] din_4_12,
    input din_valid_4_12,
    input [NF_WIDTH-1:0] din_4_13,
    input din_valid_4_13,
    input [NF_WIDTH-1:0] din_4_14,
    input din_valid_4_14,
    input [NF_WIDTH-1:0] din_4_15,
    input din_valid_4_15,
    input [NF_WIDTH-1:0] din_5_0,
    input din_valid_5_0,
    input [NF_WIDTH-1:0] din_5_1,
    input din_valid_5_1,
    input [NF_WIDTH-1:0] din_5_2,
    input din_valid_5_2,
    input [NF_WIDTH-1:0] din_5_3,
    input din_valid_5_3,
    input [NF_WIDTH-1:0] din_5_4,
    input din_valid_5_4,
    input [NF_WIDTH-1:0] din_5_5,
    input din_valid_5_5,
    input [NF_WIDTH-1:0] din_5_6,
    input din_valid_5_6,
    input [NF_WIDTH-1:0] din_5_7,
    input din_valid_5_7,
    input [NF_WIDTH-1:0] din_5_8,
    input din_valid_5_8,
    input [NF_WIDTH-1:0] din_5_9,
    input din_valid_5_9,
    input [NF_WIDTH-1:0] din_5_10,
    input din_valid_5_10,
    input [NF_WIDTH-1:0] din_5_11,
    input din_valid_5_11,
    input [NF_WIDTH-1:0] din_5_12,
    input din_valid_5_12,
    input [NF_WIDTH-1:0] din_5_13,
    input din_valid_5_13,
    input [NF_WIDTH-1:0] din_5_14,
    input din_valid_5_14,
    input [NF_WIDTH-1:0] din_5_15,
    input din_valid_5_15,
    input [NF_WIDTH-1:0] din_6_0,
    input din_valid_6_0,
    input [NF_WIDTH-1:0] din_6_1,
    input din_valid_6_1,
    input [NF_WIDTH-1:0] din_6_2,
    input din_valid_6_2,
    input [NF_WIDTH-1:0] din_6_3,
    input din_valid_6_3,
    input [NF_WIDTH-1:0] din_6_4,
    input din_valid_6_4,
    input [NF_WIDTH-1:0] din_6_5,
    input din_valid_6_5,
    input [NF_WIDTH-1:0] din_6_6,
    input din_valid_6_6,
    input [NF_WIDTH-1:0] din_6_7,
    input din_valid_6_7,
    input [NF_WIDTH-1:0] din_6_8,
    input din_valid_6_8,
    input [NF_WIDTH-1:0] din_6_9,
    input din_valid_6_9,
    input [NF_WIDTH-1:0] din_6_10,
    input din_valid_6_10,
    input [NF_WIDTH-1:0] din_6_11,
    input din_valid_6_11,
    input [NF_WIDTH-1:0] din_6_12,
    input din_valid_6_12,
    input [NF_WIDTH-1:0] din_6_13,
    input din_valid_6_13,
    input [NF_WIDTH-1:0] din_6_14,
    input din_valid_6_14,
    input [NF_WIDTH-1:0] din_6_15,
    input din_valid_6_15,
    input [NF_WIDTH-1:0] din_7_0,
    input din_valid_7_0,
    input [NF_WIDTH-1:0] din_7_1,
    input din_valid_7_1,
    input [NF_WIDTH-1:0] din_7_2,
    input din_valid_7_2,
    input [NF_WIDTH-1:0] din_7_3,
    input din_valid_7_3,
    input [NF_WIDTH-1:0] din_7_4,
    input din_valid_7_4,
    input [NF_WIDTH-1:0] din_7_5,
    input din_valid_7_5,
    input [NF_WIDTH-1:0] din_7_6,
    input din_valid_7_6,
    input [NF_WIDTH-1:0] din_7_7,
    input din_valid_7_7,
    input [NF_WIDTH-1:0] din_7_8,
    input din_valid_7_8,
    input [NF_WIDTH-1:0] din_7_9,
    input din_valid_7_9,
    input [NF_WIDTH-1:0] din_7_10,
    input din_valid_7_10,
    input [NF_WIDTH-1:0] din_7_11,
    input din_valid_7_11,
    input [NF_WIDTH-1:0] din_7_12,
    input din_valid_7_12,
    input [NF_WIDTH-1:0] din_7_13,
    input din_valid_7_13,
    input [NF_WIDTH-1:0] din_7_14,
    input din_valid_7_14,
    input [NF_WIDTH-1:0] din_7_15,
    input din_valid_7_15,
    input  last
);

//L1
logic [BUCKET_BITS-1:0] index_trunc_0_0;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_0;
logic                    l1_valid_0_0;
logic [BUCKET_BITS-1:0] index_trunc_0_1;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_1;
logic                    l1_valid_0_1;
logic [BUCKET_BITS-1:0] index_trunc_0_2;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_2;
logic                    l1_valid_0_2;
logic [BUCKET_BITS-1:0] index_trunc_0_3;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_3;
logic                    l1_valid_0_3;
logic [BUCKET_BITS-1:0] index_trunc_0_4;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_4;
logic                    l1_valid_0_4;
logic [BUCKET_BITS-1:0] index_trunc_0_5;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_5;
logic                    l1_valid_0_5;
logic [BUCKET_BITS-1:0] index_trunc_0_6;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_6;
logic                    l1_valid_0_6;
logic [BUCKET_BITS-1:0] index_trunc_0_7;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_7;
logic                    l1_valid_0_7;
logic [BUCKET_BITS-1:0] index_trunc_0_8;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_8;
logic                    l1_valid_0_8;
logic [BUCKET_BITS-1:0] index_trunc_0_9;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_9;
logic                    l1_valid_0_9;
logic [BUCKET_BITS-1:0] index_trunc_0_10;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_10;
logic                    l1_valid_0_10;
logic [BUCKET_BITS-1:0] index_trunc_0_11;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_11;
logic                    l1_valid_0_11;
logic [BUCKET_BITS-1:0] index_trunc_0_12;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_12;
logic                    l1_valid_0_12;
logic [BUCKET_BITS-1:0] index_trunc_0_13;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_13;
logic                    l1_valid_0_13;
logic [BUCKET_BITS-1:0] index_trunc_0_14;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_14;
logic                    l1_valid_0_14;
logic [BUCKET_BITS-1:0] index_trunc_0_15;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_0_15;
logic                    l1_valid_0_15;
logic [BUCKET_BITS-1:0] index_trunc_1_0;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_0;
logic                    l1_valid_1_0;
logic [BUCKET_BITS-1:0] index_trunc_1_1;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_1;
logic                    l1_valid_1_1;
logic [BUCKET_BITS-1:0] index_trunc_1_2;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_2;
logic                    l1_valid_1_2;
logic [BUCKET_BITS-1:0] index_trunc_1_3;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_3;
logic                    l1_valid_1_3;
logic [BUCKET_BITS-1:0] index_trunc_1_4;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_4;
logic                    l1_valid_1_4;
logic [BUCKET_BITS-1:0] index_trunc_1_5;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_5;
logic                    l1_valid_1_5;
logic [BUCKET_BITS-1:0] index_trunc_1_6;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_6;
logic                    l1_valid_1_6;
logic [BUCKET_BITS-1:0] index_trunc_1_7;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_7;
logic                    l1_valid_1_7;
logic [BUCKET_BITS-1:0] index_trunc_1_8;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_8;
logic                    l1_valid_1_8;
logic [BUCKET_BITS-1:0] index_trunc_1_9;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_9;
logic                    l1_valid_1_9;
logic [BUCKET_BITS-1:0] index_trunc_1_10;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_10;
logic                    l1_valid_1_10;
logic [BUCKET_BITS-1:0] index_trunc_1_11;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_11;
logic                    l1_valid_1_11;
logic [BUCKET_BITS-1:0] index_trunc_1_12;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_12;
logic                    l1_valid_1_12;
logic [BUCKET_BITS-1:0] index_trunc_1_13;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_13;
logic                    l1_valid_1_13;
logic [BUCKET_BITS-1:0] index_trunc_1_14;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_14;
logic                    l1_valid_1_14;
logic [BUCKET_BITS-1:0] index_trunc_1_15;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_1_15;
logic                    l1_valid_1_15;
logic [BUCKET_BITS-1:0] index_trunc_2_0;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_0;
logic                    l1_valid_2_0;
logic [BUCKET_BITS-1:0] index_trunc_2_1;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_1;
logic                    l1_valid_2_1;
logic [BUCKET_BITS-1:0] index_trunc_2_2;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_2;
logic                    l1_valid_2_2;
logic [BUCKET_BITS-1:0] index_trunc_2_3;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_3;
logic                    l1_valid_2_3;
logic [BUCKET_BITS-1:0] index_trunc_2_4;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_4;
logic                    l1_valid_2_4;
logic [BUCKET_BITS-1:0] index_trunc_2_5;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_5;
logic                    l1_valid_2_5;
logic [BUCKET_BITS-1:0] index_trunc_2_6;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_6;
logic                    l1_valid_2_6;
logic [BUCKET_BITS-1:0] index_trunc_2_7;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_7;
logic                    l1_valid_2_7;
logic [BUCKET_BITS-1:0] index_trunc_2_8;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_8;
logic                    l1_valid_2_8;
logic [BUCKET_BITS-1:0] index_trunc_2_9;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_9;
logic                    l1_valid_2_9;
logic [BUCKET_BITS-1:0] index_trunc_2_10;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_10;
logic                    l1_valid_2_10;
logic [BUCKET_BITS-1:0] index_trunc_2_11;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_11;
logic                    l1_valid_2_11;
logic [BUCKET_BITS-1:0] index_trunc_2_12;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_12;
logic                    l1_valid_2_12;
logic [BUCKET_BITS-1:0] index_trunc_2_13;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_13;
logic                    l1_valid_2_13;
logic [BUCKET_BITS-1:0] index_trunc_2_14;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_14;
logic                    l1_valid_2_14;
logic [BUCKET_BITS-1:0] index_trunc_2_15;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_2_15;
logic                    l1_valid_2_15;
logic [BUCKET_BITS-1:0] index_trunc_3_0;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_0;
logic                    l1_valid_3_0;
logic [BUCKET_BITS-1:0] index_trunc_3_1;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_1;
logic                    l1_valid_3_1;
logic [BUCKET_BITS-1:0] index_trunc_3_2;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_2;
logic                    l1_valid_3_2;
logic [BUCKET_BITS-1:0] index_trunc_3_3;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_3;
logic                    l1_valid_3_3;
logic [BUCKET_BITS-1:0] index_trunc_3_4;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_4;
logic                    l1_valid_3_4;
logic [BUCKET_BITS-1:0] index_trunc_3_5;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_5;
logic                    l1_valid_3_5;
logic [BUCKET_BITS-1:0] index_trunc_3_6;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_6;
logic                    l1_valid_3_6;
logic [BUCKET_BITS-1:0] index_trunc_3_7;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_7;
logic                    l1_valid_3_7;
logic [BUCKET_BITS-1:0] index_trunc_3_8;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_8;
logic                    l1_valid_3_8;
logic [BUCKET_BITS-1:0] index_trunc_3_9;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_9;
logic                    l1_valid_3_9;
logic [BUCKET_BITS-1:0] index_trunc_3_10;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_10;
logic                    l1_valid_3_10;
logic [BUCKET_BITS-1:0] index_trunc_3_11;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_11;
logic                    l1_valid_3_11;
logic [BUCKET_BITS-1:0] index_trunc_3_12;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_12;
logic                    l1_valid_3_12;
logic [BUCKET_BITS-1:0] index_trunc_3_13;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_13;
logic                    l1_valid_3_13;
logic [BUCKET_BITS-1:0] index_trunc_3_14;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_14;
logic                    l1_valid_3_14;
logic [BUCKET_BITS-1:0] index_trunc_3_15;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_3_15;
logic                    l1_valid_3_15;
logic [BUCKET_BITS-1:0] index_trunc_4_0;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_0;
logic                    l1_valid_4_0;
logic [BUCKET_BITS-1:0] index_trunc_4_1;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_1;
logic                    l1_valid_4_1;
logic [BUCKET_BITS-1:0] index_trunc_4_2;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_2;
logic                    l1_valid_4_2;
logic [BUCKET_BITS-1:0] index_trunc_4_3;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_3;
logic                    l1_valid_4_3;
logic [BUCKET_BITS-1:0] index_trunc_4_4;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_4;
logic                    l1_valid_4_4;
logic [BUCKET_BITS-1:0] index_trunc_4_5;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_5;
logic                    l1_valid_4_5;
logic [BUCKET_BITS-1:0] index_trunc_4_6;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_6;
logic                    l1_valid_4_6;
logic [BUCKET_BITS-1:0] index_trunc_4_7;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_7;
logic                    l1_valid_4_7;
logic [BUCKET_BITS-1:0] index_trunc_4_8;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_8;
logic                    l1_valid_4_8;
logic [BUCKET_BITS-1:0] index_trunc_4_9;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_9;
logic                    l1_valid_4_9;
logic [BUCKET_BITS-1:0] index_trunc_4_10;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_10;
logic                    l1_valid_4_10;
logic [BUCKET_BITS-1:0] index_trunc_4_11;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_11;
logic                    l1_valid_4_11;
logic [BUCKET_BITS-1:0] index_trunc_4_12;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_12;
logic                    l1_valid_4_12;
logic [BUCKET_BITS-1:0] index_trunc_4_13;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_13;
logic                    l1_valid_4_13;
logic [BUCKET_BITS-1:0] index_trunc_4_14;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_14;
logic                    l1_valid_4_14;
logic [BUCKET_BITS-1:0] index_trunc_4_15;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_4_15;
logic                    l1_valid_4_15;
logic [BUCKET_BITS-1:0] index_trunc_5_0;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_0;
logic                    l1_valid_5_0;
logic [BUCKET_BITS-1:0] index_trunc_5_1;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_1;
logic                    l1_valid_5_1;
logic [BUCKET_BITS-1:0] index_trunc_5_2;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_2;
logic                    l1_valid_5_2;
logic [BUCKET_BITS-1:0] index_trunc_5_3;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_3;
logic                    l1_valid_5_3;
logic [BUCKET_BITS-1:0] index_trunc_5_4;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_4;
logic                    l1_valid_5_4;
logic [BUCKET_BITS-1:0] index_trunc_5_5;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_5;
logic                    l1_valid_5_5;
logic [BUCKET_BITS-1:0] index_trunc_5_6;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_6;
logic                    l1_valid_5_6;
logic [BUCKET_BITS-1:0] index_trunc_5_7;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_7;
logic                    l1_valid_5_7;
logic [BUCKET_BITS-1:0] index_trunc_5_8;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_8;
logic                    l1_valid_5_8;
logic [BUCKET_BITS-1:0] index_trunc_5_9;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_9;
logic                    l1_valid_5_9;
logic [BUCKET_BITS-1:0] index_trunc_5_10;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_10;
logic                    l1_valid_5_10;
logic [BUCKET_BITS-1:0] index_trunc_5_11;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_11;
logic                    l1_valid_5_11;
logic [BUCKET_BITS-1:0] index_trunc_5_12;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_12;
logic                    l1_valid_5_12;
logic [BUCKET_BITS-1:0] index_trunc_5_13;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_13;
logic                    l1_valid_5_13;
logic [BUCKET_BITS-1:0] index_trunc_5_14;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_14;
logic                    l1_valid_5_14;
logic [BUCKET_BITS-1:0] index_trunc_5_15;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_5_15;
logic                    l1_valid_5_15;
logic [BUCKET_BITS-1:0] index_trunc_6_0;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_0;
logic                    l1_valid_6_0;
logic [BUCKET_BITS-1:0] index_trunc_6_1;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_1;
logic                    l1_valid_6_1;
logic [BUCKET_BITS-1:0] index_trunc_6_2;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_2;
logic                    l1_valid_6_2;
logic [BUCKET_BITS-1:0] index_trunc_6_3;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_3;
logic                    l1_valid_6_3;
logic [BUCKET_BITS-1:0] index_trunc_6_4;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_4;
logic                    l1_valid_6_4;
logic [BUCKET_BITS-1:0] index_trunc_6_5;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_5;
logic                    l1_valid_6_5;
logic [BUCKET_BITS-1:0] index_trunc_6_6;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_6;
logic                    l1_valid_6_6;
logic [BUCKET_BITS-1:0] index_trunc_6_7;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_7;
logic                    l1_valid_6_7;
logic [BUCKET_BITS-1:0] index_trunc_6_8;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_8;
logic                    l1_valid_6_8;
logic [BUCKET_BITS-1:0] index_trunc_6_9;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_9;
logic                    l1_valid_6_9;
logic [BUCKET_BITS-1:0] index_trunc_6_10;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_10;
logic                    l1_valid_6_10;
logic [BUCKET_BITS-1:0] index_trunc_6_11;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_11;
logic                    l1_valid_6_11;
logic [BUCKET_BITS-1:0] index_trunc_6_12;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_12;
logic                    l1_valid_6_12;
logic [BUCKET_BITS-1:0] index_trunc_6_13;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_13;
logic                    l1_valid_6_13;
logic [BUCKET_BITS-1:0] index_trunc_6_14;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_14;
logic                    l1_valid_6_14;
logic [BUCKET_BITS-1:0] index_trunc_6_15;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_6_15;
logic                    l1_valid_6_15;
logic [BUCKET_BITS-1:0] index_trunc_7_0;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_0;
logic                    l1_valid_7_0;
logic [BUCKET_BITS-1:0] index_trunc_7_1;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_1;
logic                    l1_valid_7_1;
logic [BUCKET_BITS-1:0] index_trunc_7_2;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_2;
logic                    l1_valid_7_2;
logic [BUCKET_BITS-1:0] index_trunc_7_3;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_3;
logic                    l1_valid_7_3;
logic [BUCKET_BITS-1:0] index_trunc_7_4;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_4;
logic                    l1_valid_7_4;
logic [BUCKET_BITS-1:0] index_trunc_7_5;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_5;
logic                    l1_valid_7_5;
logic [BUCKET_BITS-1:0] index_trunc_7_6;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_6;
logic                    l1_valid_7_6;
logic [BUCKET_BITS-1:0] index_trunc_7_7;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_7;
logic                    l1_valid_7_7;
logic [BUCKET_BITS-1:0] index_trunc_7_8;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_8;
logic                    l1_valid_7_8;
logic [BUCKET_BITS-1:0] index_trunc_7_9;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_9;
logic                    l1_valid_7_9;
logic [BUCKET_BITS-1:0] index_trunc_7_10;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_10;
logic                    l1_valid_7_10;
logic [BUCKET_BITS-1:0] index_trunc_7_11;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_11;
logic                    l1_valid_7_11;
logic [BUCKET_BITS-1:0] index_trunc_7_12;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_12;
logic                    l1_valid_7_12;
logic [BUCKET_BITS-1:0] index_trunc_7_13;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_13;
logic                    l1_valid_7_13;
logic [BUCKET_BITS-1:0] index_trunc_7_14;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_14;
logic                    l1_valid_7_14;
logic [BUCKET_BITS-1:0] index_trunc_7_15;
logic [BUCKET_WIDTH-1:0] l1_sub_fp_7_15;
logic                    l1_valid_7_15;

//L2
logic [BUCKET_WIDTH-1:0] l2_sub_fp_0_0;
logic                    l2_valid_0_0;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_0_1;
logic                    l2_valid_0_1;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_0_2;
logic                    l2_valid_0_2;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_0_3;
logic                    l2_valid_0_3;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_0_4;
logic                    l2_valid_0_4;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_0_5;
logic                    l2_valid_0_5;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_0_6;
logic                    l2_valid_0_6;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_0_7;
logic                    l2_valid_0_7;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_1_0;
logic                    l2_valid_1_0;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_1_1;
logic                    l2_valid_1_1;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_1_2;
logic                    l2_valid_1_2;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_1_3;
logic                    l2_valid_1_3;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_1_4;
logic                    l2_valid_1_4;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_1_5;
logic                    l2_valid_1_5;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_1_6;
logic                    l2_valid_1_6;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_1_7;
logic                    l2_valid_1_7;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_2_0;
logic                    l2_valid_2_0;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_2_1;
logic                    l2_valid_2_1;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_2_2;
logic                    l2_valid_2_2;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_2_3;
logic                    l2_valid_2_3;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_2_4;
logic                    l2_valid_2_4;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_2_5;
logic                    l2_valid_2_5;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_2_6;
logic                    l2_valid_2_6;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_2_7;
logic                    l2_valid_2_7;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_3_0;
logic                    l2_valid_3_0;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_3_1;
logic                    l2_valid_3_1;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_3_2;
logic                    l2_valid_3_2;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_3_3;
logic                    l2_valid_3_3;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_3_4;
logic                    l2_valid_3_4;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_3_5;
logic                    l2_valid_3_5;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_3_6;
logic                    l2_valid_3_6;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_3_7;
logic                    l2_valid_3_7;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_4_0;
logic                    l2_valid_4_0;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_4_1;
logic                    l2_valid_4_1;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_4_2;
logic                    l2_valid_4_2;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_4_3;
logic                    l2_valid_4_3;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_4_4;
logic                    l2_valid_4_4;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_4_5;
logic                    l2_valid_4_5;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_4_6;
logic                    l2_valid_4_6;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_4_7;
logic                    l2_valid_4_7;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_5_0;
logic                    l2_valid_5_0;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_5_1;
logic                    l2_valid_5_1;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_5_2;
logic                    l2_valid_5_2;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_5_3;
logic                    l2_valid_5_3;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_5_4;
logic                    l2_valid_5_4;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_5_5;
logic                    l2_valid_5_5;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_5_6;
logic                    l2_valid_5_6;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_5_7;
logic                    l2_valid_5_7;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_6_0;
logic                    l2_valid_6_0;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_6_1;
logic                    l2_valid_6_1;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_6_2;
logic                    l2_valid_6_2;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_6_3;
logic                    l2_valid_6_3;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_6_4;
logic                    l2_valid_6_4;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_6_5;
logic                    l2_valid_6_5;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_6_6;
logic                    l2_valid_6_6;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_6_7;
logic                    l2_valid_6_7;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_7_0;
logic                    l2_valid_7_0;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_7_1;
logic                    l2_valid_7_1;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_7_2;
logic                    l2_valid_7_2;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_7_3;
logic                    l2_valid_7_3;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_7_4;
logic                    l2_valid_7_4;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_7_5;
logic                    l2_valid_7_5;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_7_6;
logic                    l2_valid_7_6;
logic [BUCKET_WIDTH-1:0] l2_sub_fp_7_7;
logic                    l2_valid_7_7;

//L3
logic [BUCKET_WIDTH-1:0] l3_sub_fp_0_0;
logic                    l3_valid_0_0;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_0_1;
logic                    l3_valid_0_1;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_0_2;
logic                    l3_valid_0_2;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_0_3;
logic                    l3_valid_0_3;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_1_0;
logic                    l3_valid_1_0;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_1_1;
logic                    l3_valid_1_1;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_1_2;
logic                    l3_valid_1_2;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_1_3;
logic                    l3_valid_1_3;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_2_0;
logic                    l3_valid_2_0;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_2_1;
logic                    l3_valid_2_1;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_2_2;
logic                    l3_valid_2_2;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_2_3;
logic                    l3_valid_2_3;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_3_0;
logic                    l3_valid_3_0;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_3_1;
logic                    l3_valid_3_1;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_3_2;
logic                    l3_valid_3_2;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_3_3;
logic                    l3_valid_3_3;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_4_0;
logic                    l3_valid_4_0;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_4_1;
logic                    l3_valid_4_1;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_4_2;
logic                    l3_valid_4_2;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_4_3;
logic                    l3_valid_4_3;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_5_0;
logic                    l3_valid_5_0;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_5_1;
logic                    l3_valid_5_1;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_5_2;
logic                    l3_valid_5_2;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_5_3;
logic                    l3_valid_5_3;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_6_0;
logic                    l3_valid_6_0;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_6_1;
logic                    l3_valid_6_1;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_6_2;
logic                    l3_valid_6_2;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_6_3;
logic                    l3_valid_6_3;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_7_0;
logic                    l3_valid_7_0;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_7_1;
logic                    l3_valid_7_1;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_7_2;
logic                    l3_valid_7_2;
logic [BUCKET_WIDTH-1:0] l3_sub_fp_7_3;
logic                    l3_valid_7_3;

//L4
logic [BUCKET_WIDTH-1:0] l4_sub_fp_0;
logic                    l4_valid_0;
logic [BUCKET_WIDTH-1:0] l4_sub_fp_1;
logic                    l4_valid_1;
logic [BUCKET_WIDTH-1:0] l4_sub_fp_2;
logic                    l4_valid_2;
logic [BUCKET_WIDTH-1:0] l4_sub_fp_3;
logic                    l4_valid_3;
logic [BUCKET_WIDTH-1:0] l4_sub_fp_4;
logic                    l4_valid_4;
logic [BUCKET_WIDTH-1:0] l4_sub_fp_5;
logic                    l4_valid_5;
logic [BUCKET_WIDTH-1:0] l4_sub_fp_6;
logic                    l4_valid_6;
logic [BUCKET_WIDTH-1:0] l4_sub_fp_7;
logic                    l4_valid_7;

//L5
logic [BUCKET_WIDTH-1:0] sub_fp_0;
logic [BUCKET_WIDTH-1:0] sub_fp_1;
logic [BUCKET_WIDTH-1:0] sub_fp_2;
logic [BUCKET_WIDTH-1:0] sub_fp_3;
logic [BUCKET_WIDTH-1:0] sub_fp_4;
logic [BUCKET_WIDTH-1:0] sub_fp_5;
logic [BUCKET_WIDTH-1:0] sub_fp_6;
logic [BUCKET_WIDTH-1:0] sub_fp_7;

logic last_r1;
logic last_r2;
logic last_r3;
logic last_r4;

assign index_trunc_0_0 = din_0_0[BUCKET_BITS-1:0];
assign index_trunc_0_1 = din_0_1[BUCKET_BITS-1:0];
assign index_trunc_0_2 = din_0_2[BUCKET_BITS-1:0];
assign index_trunc_0_3 = din_0_3[BUCKET_BITS-1:0];
assign index_trunc_0_4 = din_0_4[BUCKET_BITS-1:0];
assign index_trunc_0_5 = din_0_5[BUCKET_BITS-1:0];
assign index_trunc_0_6 = din_0_6[BUCKET_BITS-1:0];
assign index_trunc_0_7 = din_0_7[BUCKET_BITS-1:0];
assign index_trunc_0_8 = din_0_8[BUCKET_BITS-1:0];
assign index_trunc_0_9 = din_0_9[BUCKET_BITS-1:0];
assign index_trunc_0_10 = din_0_10[BUCKET_BITS-1:0];
assign index_trunc_0_11 = din_0_11[BUCKET_BITS-1:0];
assign index_trunc_0_12 = din_0_12[BUCKET_BITS-1:0];
assign index_trunc_0_13 = din_0_13[BUCKET_BITS-1:0];
assign index_trunc_0_14 = din_0_14[BUCKET_BITS-1:0];
assign index_trunc_0_15 = din_0_15[BUCKET_BITS-1:0];
assign index_trunc_1_0 = din_1_0[BUCKET_BITS-1:0];
assign index_trunc_1_1 = din_1_1[BUCKET_BITS-1:0];
assign index_trunc_1_2 = din_1_2[BUCKET_BITS-1:0];
assign index_trunc_1_3 = din_1_3[BUCKET_BITS-1:0];
assign index_trunc_1_4 = din_1_4[BUCKET_BITS-1:0];
assign index_trunc_1_5 = din_1_5[BUCKET_BITS-1:0];
assign index_trunc_1_6 = din_1_6[BUCKET_BITS-1:0];
assign index_trunc_1_7 = din_1_7[BUCKET_BITS-1:0];
assign index_trunc_1_8 = din_1_8[BUCKET_BITS-1:0];
assign index_trunc_1_9 = din_1_9[BUCKET_BITS-1:0];
assign index_trunc_1_10 = din_1_10[BUCKET_BITS-1:0];
assign index_trunc_1_11 = din_1_11[BUCKET_BITS-1:0];
assign index_trunc_1_12 = din_1_12[BUCKET_BITS-1:0];
assign index_trunc_1_13 = din_1_13[BUCKET_BITS-1:0];
assign index_trunc_1_14 = din_1_14[BUCKET_BITS-1:0];
assign index_trunc_1_15 = din_1_15[BUCKET_BITS-1:0];
assign index_trunc_2_0 = din_2_0[BUCKET_BITS-1:0];
assign index_trunc_2_1 = din_2_1[BUCKET_BITS-1:0];
assign index_trunc_2_2 = din_2_2[BUCKET_BITS-1:0];
assign index_trunc_2_3 = din_2_3[BUCKET_BITS-1:0];
assign index_trunc_2_4 = din_2_4[BUCKET_BITS-1:0];
assign index_trunc_2_5 = din_2_5[BUCKET_BITS-1:0];
assign index_trunc_2_6 = din_2_6[BUCKET_BITS-1:0];
assign index_trunc_2_7 = din_2_7[BUCKET_BITS-1:0];
assign index_trunc_2_8 = din_2_8[BUCKET_BITS-1:0];
assign index_trunc_2_9 = din_2_9[BUCKET_BITS-1:0];
assign index_trunc_2_10 = din_2_10[BUCKET_BITS-1:0];
assign index_trunc_2_11 = din_2_11[BUCKET_BITS-1:0];
assign index_trunc_2_12 = din_2_12[BUCKET_BITS-1:0];
assign index_trunc_2_13 = din_2_13[BUCKET_BITS-1:0];
assign index_trunc_2_14 = din_2_14[BUCKET_BITS-1:0];
assign index_trunc_2_15 = din_2_15[BUCKET_BITS-1:0];
assign index_trunc_3_0 = din_3_0[BUCKET_BITS-1:0];
assign index_trunc_3_1 = din_3_1[BUCKET_BITS-1:0];
assign index_trunc_3_2 = din_3_2[BUCKET_BITS-1:0];
assign index_trunc_3_3 = din_3_3[BUCKET_BITS-1:0];
assign index_trunc_3_4 = din_3_4[BUCKET_BITS-1:0];
assign index_trunc_3_5 = din_3_5[BUCKET_BITS-1:0];
assign index_trunc_3_6 = din_3_6[BUCKET_BITS-1:0];
assign index_trunc_3_7 = din_3_7[BUCKET_BITS-1:0];
assign index_trunc_3_8 = din_3_8[BUCKET_BITS-1:0];
assign index_trunc_3_9 = din_3_9[BUCKET_BITS-1:0];
assign index_trunc_3_10 = din_3_10[BUCKET_BITS-1:0];
assign index_trunc_3_11 = din_3_11[BUCKET_BITS-1:0];
assign index_trunc_3_12 = din_3_12[BUCKET_BITS-1:0];
assign index_trunc_3_13 = din_3_13[BUCKET_BITS-1:0];
assign index_trunc_3_14 = din_3_14[BUCKET_BITS-1:0];
assign index_trunc_3_15 = din_3_15[BUCKET_BITS-1:0];
assign index_trunc_4_0 = din_4_0[BUCKET_BITS-1:0];
assign index_trunc_4_1 = din_4_1[BUCKET_BITS-1:0];
assign index_trunc_4_2 = din_4_2[BUCKET_BITS-1:0];
assign index_trunc_4_3 = din_4_3[BUCKET_BITS-1:0];
assign index_trunc_4_4 = din_4_4[BUCKET_BITS-1:0];
assign index_trunc_4_5 = din_4_5[BUCKET_BITS-1:0];
assign index_trunc_4_6 = din_4_6[BUCKET_BITS-1:0];
assign index_trunc_4_7 = din_4_7[BUCKET_BITS-1:0];
assign index_trunc_4_8 = din_4_8[BUCKET_BITS-1:0];
assign index_trunc_4_9 = din_4_9[BUCKET_BITS-1:0];
assign index_trunc_4_10 = din_4_10[BUCKET_BITS-1:0];
assign index_trunc_4_11 = din_4_11[BUCKET_BITS-1:0];
assign index_trunc_4_12 = din_4_12[BUCKET_BITS-1:0];
assign index_trunc_4_13 = din_4_13[BUCKET_BITS-1:0];
assign index_trunc_4_14 = din_4_14[BUCKET_BITS-1:0];
assign index_trunc_4_15 = din_4_15[BUCKET_BITS-1:0];
assign index_trunc_5_0 = din_5_0[BUCKET_BITS-1:0];
assign index_trunc_5_1 = din_5_1[BUCKET_BITS-1:0];
assign index_trunc_5_2 = din_5_2[BUCKET_BITS-1:0];
assign index_trunc_5_3 = din_5_3[BUCKET_BITS-1:0];
assign index_trunc_5_4 = din_5_4[BUCKET_BITS-1:0];
assign index_trunc_5_5 = din_5_5[BUCKET_BITS-1:0];
assign index_trunc_5_6 = din_5_6[BUCKET_BITS-1:0];
assign index_trunc_5_7 = din_5_7[BUCKET_BITS-1:0];
assign index_trunc_5_8 = din_5_8[BUCKET_BITS-1:0];
assign index_trunc_5_9 = din_5_9[BUCKET_BITS-1:0];
assign index_trunc_5_10 = din_5_10[BUCKET_BITS-1:0];
assign index_trunc_5_11 = din_5_11[BUCKET_BITS-1:0];
assign index_trunc_5_12 = din_5_12[BUCKET_BITS-1:0];
assign index_trunc_5_13 = din_5_13[BUCKET_BITS-1:0];
assign index_trunc_5_14 = din_5_14[BUCKET_BITS-1:0];
assign index_trunc_5_15 = din_5_15[BUCKET_BITS-1:0];
assign index_trunc_6_0 = din_6_0[BUCKET_BITS-1:0];
assign index_trunc_6_1 = din_6_1[BUCKET_BITS-1:0];
assign index_trunc_6_2 = din_6_2[BUCKET_BITS-1:0];
assign index_trunc_6_3 = din_6_3[BUCKET_BITS-1:0];
assign index_trunc_6_4 = din_6_4[BUCKET_BITS-1:0];
assign index_trunc_6_5 = din_6_5[BUCKET_BITS-1:0];
assign index_trunc_6_6 = din_6_6[BUCKET_BITS-1:0];
assign index_trunc_6_7 = din_6_7[BUCKET_BITS-1:0];
assign index_trunc_6_8 = din_6_8[BUCKET_BITS-1:0];
assign index_trunc_6_9 = din_6_9[BUCKET_BITS-1:0];
assign index_trunc_6_10 = din_6_10[BUCKET_BITS-1:0];
assign index_trunc_6_11 = din_6_11[BUCKET_BITS-1:0];
assign index_trunc_6_12 = din_6_12[BUCKET_BITS-1:0];
assign index_trunc_6_13 = din_6_13[BUCKET_BITS-1:0];
assign index_trunc_6_14 = din_6_14[BUCKET_BITS-1:0];
assign index_trunc_6_15 = din_6_15[BUCKET_BITS-1:0];
assign index_trunc_7_0 = din_7_0[BUCKET_BITS-1:0];
assign index_trunc_7_1 = din_7_1[BUCKET_BITS-1:0];
assign index_trunc_7_2 = din_7_2[BUCKET_BITS-1:0];
assign index_trunc_7_3 = din_7_3[BUCKET_BITS-1:0];
assign index_trunc_7_4 = din_7_4[BUCKET_BITS-1:0];
assign index_trunc_7_5 = din_7_5[BUCKET_BITS-1:0];
assign index_trunc_7_6 = din_7_6[BUCKET_BITS-1:0];
assign index_trunc_7_7 = din_7_7[BUCKET_BITS-1:0];
assign index_trunc_7_8 = din_7_8[BUCKET_BITS-1:0];
assign index_trunc_7_9 = din_7_9[BUCKET_BITS-1:0];
assign index_trunc_7_10 = din_7_10[BUCKET_BITS-1:0];
assign index_trunc_7_11 = din_7_11[BUCKET_BITS-1:0];
assign index_trunc_7_12 = din_7_12[BUCKET_BITS-1:0];
assign index_trunc_7_13 = din_7_13[BUCKET_BITS-1:0];
assign index_trunc_7_14 = din_7_14[BUCKET_BITS-1:0];
assign index_trunc_7_15 = din_7_15[BUCKET_BITS-1:0];


//Layer 1
always@(posedge clk)begin
    l1_sub_fp_0_0 <= 0;
    l1_valid_0_0 <= 0;
    if(din_valid_0_0)begin
        l1_sub_fp_0_0 <= 1 << index_trunc_0_0;
        l1_valid_0_0 <= 1;
    end
    l1_sub_fp_0_1 <= 0;
    l1_valid_0_1 <= 0;
    if(din_valid_0_1)begin
        l1_sub_fp_0_1 <= 1 << index_trunc_0_1;
        l1_valid_0_1 <= 1;
    end
    l1_sub_fp_0_2 <= 0;
    l1_valid_0_2 <= 0;
    if(din_valid_0_2)begin
        l1_sub_fp_0_2 <= 1 << index_trunc_0_2;
        l1_valid_0_2 <= 1;
    end
    l1_sub_fp_0_3 <= 0;
    l1_valid_0_3 <= 0;
    if(din_valid_0_3)begin
        l1_sub_fp_0_3 <= 1 << index_trunc_0_3;
        l1_valid_0_3 <= 1;
    end
    l1_sub_fp_0_4 <= 0;
    l1_valid_0_4 <= 0;
    if(din_valid_0_4)begin
        l1_sub_fp_0_4 <= 1 << index_trunc_0_4;
        l1_valid_0_4 <= 1;
    end
    l1_sub_fp_0_5 <= 0;
    l1_valid_0_5 <= 0;
    if(din_valid_0_5)begin
        l1_sub_fp_0_5 <= 1 << index_trunc_0_5;
        l1_valid_0_5 <= 1;
    end
    l1_sub_fp_0_6 <= 0;
    l1_valid_0_6 <= 0;
    if(din_valid_0_6)begin
        l1_sub_fp_0_6 <= 1 << index_trunc_0_6;
        l1_valid_0_6 <= 1;
    end
    l1_sub_fp_0_7 <= 0;
    l1_valid_0_7 <= 0;
    if(din_valid_0_7)begin
        l1_sub_fp_0_7 <= 1 << index_trunc_0_7;
        l1_valid_0_7 <= 1;
    end
    l1_sub_fp_0_8 <= 0;
    l1_valid_0_8 <= 0;
    if(din_valid_0_8)begin
        l1_sub_fp_0_8 <= 1 << index_trunc_0_8;
        l1_valid_0_8 <= 1;
    end
    l1_sub_fp_0_9 <= 0;
    l1_valid_0_9 <= 0;
    if(din_valid_0_9)begin
        l1_sub_fp_0_9 <= 1 << index_trunc_0_9;
        l1_valid_0_9 <= 1;
    end
    l1_sub_fp_0_10 <= 0;
    l1_valid_0_10 <= 0;
    if(din_valid_0_10)begin
        l1_sub_fp_0_10 <= 1 << index_trunc_0_10;
        l1_valid_0_10 <= 1;
    end
    l1_sub_fp_0_11 <= 0;
    l1_valid_0_11 <= 0;
    if(din_valid_0_11)begin
        l1_sub_fp_0_11 <= 1 << index_trunc_0_11;
        l1_valid_0_11 <= 1;
    end
    l1_sub_fp_0_12 <= 0;
    l1_valid_0_12 <= 0;
    if(din_valid_0_12)begin
        l1_sub_fp_0_12 <= 1 << index_trunc_0_12;
        l1_valid_0_12 <= 1;
    end
    l1_sub_fp_0_13 <= 0;
    l1_valid_0_13 <= 0;
    if(din_valid_0_13)begin
        l1_sub_fp_0_13 <= 1 << index_trunc_0_13;
        l1_valid_0_13 <= 1;
    end
    l1_sub_fp_0_14 <= 0;
    l1_valid_0_14 <= 0;
    if(din_valid_0_14)begin
        l1_sub_fp_0_14 <= 1 << index_trunc_0_14;
        l1_valid_0_14 <= 1;
    end
    l1_sub_fp_0_15 <= 0;
    l1_valid_0_15 <= 0;
    if(din_valid_0_15)begin
        l1_sub_fp_0_15 <= 1 << index_trunc_0_15;
        l1_valid_0_15 <= 1;
    end
    l1_sub_fp_1_0 <= 0;
    l1_valid_1_0 <= 0;
    if(din_valid_1_0)begin
        l1_sub_fp_1_0 <= 1 << index_trunc_1_0;
        l1_valid_1_0 <= 1;
    end
    l1_sub_fp_1_1 <= 0;
    l1_valid_1_1 <= 0;
    if(din_valid_1_1)begin
        l1_sub_fp_1_1 <= 1 << index_trunc_1_1;
        l1_valid_1_1 <= 1;
    end
    l1_sub_fp_1_2 <= 0;
    l1_valid_1_2 <= 0;
    if(din_valid_1_2)begin
        l1_sub_fp_1_2 <= 1 << index_trunc_1_2;
        l1_valid_1_2 <= 1;
    end
    l1_sub_fp_1_3 <= 0;
    l1_valid_1_3 <= 0;
    if(din_valid_1_3)begin
        l1_sub_fp_1_3 <= 1 << index_trunc_1_3;
        l1_valid_1_3 <= 1;
    end
    l1_sub_fp_1_4 <= 0;
    l1_valid_1_4 <= 0;
    if(din_valid_1_4)begin
        l1_sub_fp_1_4 <= 1 << index_trunc_1_4;
        l1_valid_1_4 <= 1;
    end
    l1_sub_fp_1_5 <= 0;
    l1_valid_1_5 <= 0;
    if(din_valid_1_5)begin
        l1_sub_fp_1_5 <= 1 << index_trunc_1_5;
        l1_valid_1_5 <= 1;
    end
    l1_sub_fp_1_6 <= 0;
    l1_valid_1_6 <= 0;
    if(din_valid_1_6)begin
        l1_sub_fp_1_6 <= 1 << index_trunc_1_6;
        l1_valid_1_6 <= 1;
    end
    l1_sub_fp_1_7 <= 0;
    l1_valid_1_7 <= 0;
    if(din_valid_1_7)begin
        l1_sub_fp_1_7 <= 1 << index_trunc_1_7;
        l1_valid_1_7 <= 1;
    end
    l1_sub_fp_1_8 <= 0;
    l1_valid_1_8 <= 0;
    if(din_valid_1_8)begin
        l1_sub_fp_1_8 <= 1 << index_trunc_1_8;
        l1_valid_1_8 <= 1;
    end
    l1_sub_fp_1_9 <= 0;
    l1_valid_1_9 <= 0;
    if(din_valid_1_9)begin
        l1_sub_fp_1_9 <= 1 << index_trunc_1_9;
        l1_valid_1_9 <= 1;
    end
    l1_sub_fp_1_10 <= 0;
    l1_valid_1_10 <= 0;
    if(din_valid_1_10)begin
        l1_sub_fp_1_10 <= 1 << index_trunc_1_10;
        l1_valid_1_10 <= 1;
    end
    l1_sub_fp_1_11 <= 0;
    l1_valid_1_11 <= 0;
    if(din_valid_1_11)begin
        l1_sub_fp_1_11 <= 1 << index_trunc_1_11;
        l1_valid_1_11 <= 1;
    end
    l1_sub_fp_1_12 <= 0;
    l1_valid_1_12 <= 0;
    if(din_valid_1_12)begin
        l1_sub_fp_1_12 <= 1 << index_trunc_1_12;
        l1_valid_1_12 <= 1;
    end
    l1_sub_fp_1_13 <= 0;
    l1_valid_1_13 <= 0;
    if(din_valid_1_13)begin
        l1_sub_fp_1_13 <= 1 << index_trunc_1_13;
        l1_valid_1_13 <= 1;
    end
    l1_sub_fp_1_14 <= 0;
    l1_valid_1_14 <= 0;
    if(din_valid_1_14)begin
        l1_sub_fp_1_14 <= 1 << index_trunc_1_14;
        l1_valid_1_14 <= 1;
    end
    l1_sub_fp_1_15 <= 0;
    l1_valid_1_15 <= 0;
    if(din_valid_1_15)begin
        l1_sub_fp_1_15 <= 1 << index_trunc_1_15;
        l1_valid_1_15 <= 1;
    end
    l1_sub_fp_2_0 <= 0;
    l1_valid_2_0 <= 0;
    if(din_valid_2_0)begin
        l1_sub_fp_2_0 <= 1 << index_trunc_2_0;
        l1_valid_2_0 <= 1;
    end
    l1_sub_fp_2_1 <= 0;
    l1_valid_2_1 <= 0;
    if(din_valid_2_1)begin
        l1_sub_fp_2_1 <= 1 << index_trunc_2_1;
        l1_valid_2_1 <= 1;
    end
    l1_sub_fp_2_2 <= 0;
    l1_valid_2_2 <= 0;
    if(din_valid_2_2)begin
        l1_sub_fp_2_2 <= 1 << index_trunc_2_2;
        l1_valid_2_2 <= 1;
    end
    l1_sub_fp_2_3 <= 0;
    l1_valid_2_3 <= 0;
    if(din_valid_2_3)begin
        l1_sub_fp_2_3 <= 1 << index_trunc_2_3;
        l1_valid_2_3 <= 1;
    end
    l1_sub_fp_2_4 <= 0;
    l1_valid_2_4 <= 0;
    if(din_valid_2_4)begin
        l1_sub_fp_2_4 <= 1 << index_trunc_2_4;
        l1_valid_2_4 <= 1;
    end
    l1_sub_fp_2_5 <= 0;
    l1_valid_2_5 <= 0;
    if(din_valid_2_5)begin
        l1_sub_fp_2_5 <= 1 << index_trunc_2_5;
        l1_valid_2_5 <= 1;
    end
    l1_sub_fp_2_6 <= 0;
    l1_valid_2_6 <= 0;
    if(din_valid_2_6)begin
        l1_sub_fp_2_6 <= 1 << index_trunc_2_6;
        l1_valid_2_6 <= 1;
    end
    l1_sub_fp_2_7 <= 0;
    l1_valid_2_7 <= 0;
    if(din_valid_2_7)begin
        l1_sub_fp_2_7 <= 1 << index_trunc_2_7;
        l1_valid_2_7 <= 1;
    end
    l1_sub_fp_2_8 <= 0;
    l1_valid_2_8 <= 0;
    if(din_valid_2_8)begin
        l1_sub_fp_2_8 <= 1 << index_trunc_2_8;
        l1_valid_2_8 <= 1;
    end
    l1_sub_fp_2_9 <= 0;
    l1_valid_2_9 <= 0;
    if(din_valid_2_9)begin
        l1_sub_fp_2_9 <= 1 << index_trunc_2_9;
        l1_valid_2_9 <= 1;
    end
    l1_sub_fp_2_10 <= 0;
    l1_valid_2_10 <= 0;
    if(din_valid_2_10)begin
        l1_sub_fp_2_10 <= 1 << index_trunc_2_10;
        l1_valid_2_10 <= 1;
    end
    l1_sub_fp_2_11 <= 0;
    l1_valid_2_11 <= 0;
    if(din_valid_2_11)begin
        l1_sub_fp_2_11 <= 1 << index_trunc_2_11;
        l1_valid_2_11 <= 1;
    end
    l1_sub_fp_2_12 <= 0;
    l1_valid_2_12 <= 0;
    if(din_valid_2_12)begin
        l1_sub_fp_2_12 <= 1 << index_trunc_2_12;
        l1_valid_2_12 <= 1;
    end
    l1_sub_fp_2_13 <= 0;
    l1_valid_2_13 <= 0;
    if(din_valid_2_13)begin
        l1_sub_fp_2_13 <= 1 << index_trunc_2_13;
        l1_valid_2_13 <= 1;
    end
    l1_sub_fp_2_14 <= 0;
    l1_valid_2_14 <= 0;
    if(din_valid_2_14)begin
        l1_sub_fp_2_14 <= 1 << index_trunc_2_14;
        l1_valid_2_14 <= 1;
    end
    l1_sub_fp_2_15 <= 0;
    l1_valid_2_15 <= 0;
    if(din_valid_2_15)begin
        l1_sub_fp_2_15 <= 1 << index_trunc_2_15;
        l1_valid_2_15 <= 1;
    end
    l1_sub_fp_3_0 <= 0;
    l1_valid_3_0 <= 0;
    if(din_valid_3_0)begin
        l1_sub_fp_3_0 <= 1 << index_trunc_3_0;
        l1_valid_3_0 <= 1;
    end
    l1_sub_fp_3_1 <= 0;
    l1_valid_3_1 <= 0;
    if(din_valid_3_1)begin
        l1_sub_fp_3_1 <= 1 << index_trunc_3_1;
        l1_valid_3_1 <= 1;
    end
    l1_sub_fp_3_2 <= 0;
    l1_valid_3_2 <= 0;
    if(din_valid_3_2)begin
        l1_sub_fp_3_2 <= 1 << index_trunc_3_2;
        l1_valid_3_2 <= 1;
    end
    l1_sub_fp_3_3 <= 0;
    l1_valid_3_3 <= 0;
    if(din_valid_3_3)begin
        l1_sub_fp_3_3 <= 1 << index_trunc_3_3;
        l1_valid_3_3 <= 1;
    end
    l1_sub_fp_3_4 <= 0;
    l1_valid_3_4 <= 0;
    if(din_valid_3_4)begin
        l1_sub_fp_3_4 <= 1 << index_trunc_3_4;
        l1_valid_3_4 <= 1;
    end
    l1_sub_fp_3_5 <= 0;
    l1_valid_3_5 <= 0;
    if(din_valid_3_5)begin
        l1_sub_fp_3_5 <= 1 << index_trunc_3_5;
        l1_valid_3_5 <= 1;
    end
    l1_sub_fp_3_6 <= 0;
    l1_valid_3_6 <= 0;
    if(din_valid_3_6)begin
        l1_sub_fp_3_6 <= 1 << index_trunc_3_6;
        l1_valid_3_6 <= 1;
    end
    l1_sub_fp_3_7 <= 0;
    l1_valid_3_7 <= 0;
    if(din_valid_3_7)begin
        l1_sub_fp_3_7 <= 1 << index_trunc_3_7;
        l1_valid_3_7 <= 1;
    end
    l1_sub_fp_3_8 <= 0;
    l1_valid_3_8 <= 0;
    if(din_valid_3_8)begin
        l1_sub_fp_3_8 <= 1 << index_trunc_3_8;
        l1_valid_3_8 <= 1;
    end
    l1_sub_fp_3_9 <= 0;
    l1_valid_3_9 <= 0;
    if(din_valid_3_9)begin
        l1_sub_fp_3_9 <= 1 << index_trunc_3_9;
        l1_valid_3_9 <= 1;
    end
    l1_sub_fp_3_10 <= 0;
    l1_valid_3_10 <= 0;
    if(din_valid_3_10)begin
        l1_sub_fp_3_10 <= 1 << index_trunc_3_10;
        l1_valid_3_10 <= 1;
    end
    l1_sub_fp_3_11 <= 0;
    l1_valid_3_11 <= 0;
    if(din_valid_3_11)begin
        l1_sub_fp_3_11 <= 1 << index_trunc_3_11;
        l1_valid_3_11 <= 1;
    end
    l1_sub_fp_3_12 <= 0;
    l1_valid_3_12 <= 0;
    if(din_valid_3_12)begin
        l1_sub_fp_3_12 <= 1 << index_trunc_3_12;
        l1_valid_3_12 <= 1;
    end
    l1_sub_fp_3_13 <= 0;
    l1_valid_3_13 <= 0;
    if(din_valid_3_13)begin
        l1_sub_fp_3_13 <= 1 << index_trunc_3_13;
        l1_valid_3_13 <= 1;
    end
    l1_sub_fp_3_14 <= 0;
    l1_valid_3_14 <= 0;
    if(din_valid_3_14)begin
        l1_sub_fp_3_14 <= 1 << index_trunc_3_14;
        l1_valid_3_14 <= 1;
    end
    l1_sub_fp_3_15 <= 0;
    l1_valid_3_15 <= 0;
    if(din_valid_3_15)begin
        l1_sub_fp_3_15 <= 1 << index_trunc_3_15;
        l1_valid_3_15 <= 1;
    end
    l1_sub_fp_4_0 <= 0;
    l1_valid_4_0 <= 0;
    if(din_valid_4_0)begin
        l1_sub_fp_4_0 <= 1 << index_trunc_4_0;
        l1_valid_4_0 <= 1;
    end
    l1_sub_fp_4_1 <= 0;
    l1_valid_4_1 <= 0;
    if(din_valid_4_1)begin
        l1_sub_fp_4_1 <= 1 << index_trunc_4_1;
        l1_valid_4_1 <= 1;
    end
    l1_sub_fp_4_2 <= 0;
    l1_valid_4_2 <= 0;
    if(din_valid_4_2)begin
        l1_sub_fp_4_2 <= 1 << index_trunc_4_2;
        l1_valid_4_2 <= 1;
    end
    l1_sub_fp_4_3 <= 0;
    l1_valid_4_3 <= 0;
    if(din_valid_4_3)begin
        l1_sub_fp_4_3 <= 1 << index_trunc_4_3;
        l1_valid_4_3 <= 1;
    end
    l1_sub_fp_4_4 <= 0;
    l1_valid_4_4 <= 0;
    if(din_valid_4_4)begin
        l1_sub_fp_4_4 <= 1 << index_trunc_4_4;
        l1_valid_4_4 <= 1;
    end
    l1_sub_fp_4_5 <= 0;
    l1_valid_4_5 <= 0;
    if(din_valid_4_5)begin
        l1_sub_fp_4_5 <= 1 << index_trunc_4_5;
        l1_valid_4_5 <= 1;
    end
    l1_sub_fp_4_6 <= 0;
    l1_valid_4_6 <= 0;
    if(din_valid_4_6)begin
        l1_sub_fp_4_6 <= 1 << index_trunc_4_6;
        l1_valid_4_6 <= 1;
    end
    l1_sub_fp_4_7 <= 0;
    l1_valid_4_7 <= 0;
    if(din_valid_4_7)begin
        l1_sub_fp_4_7 <= 1 << index_trunc_4_7;
        l1_valid_4_7 <= 1;
    end
    l1_sub_fp_4_8 <= 0;
    l1_valid_4_8 <= 0;
    if(din_valid_4_8)begin
        l1_sub_fp_4_8 <= 1 << index_trunc_4_8;
        l1_valid_4_8 <= 1;
    end
    l1_sub_fp_4_9 <= 0;
    l1_valid_4_9 <= 0;
    if(din_valid_4_9)begin
        l1_sub_fp_4_9 <= 1 << index_trunc_4_9;
        l1_valid_4_9 <= 1;
    end
    l1_sub_fp_4_10 <= 0;
    l1_valid_4_10 <= 0;
    if(din_valid_4_10)begin
        l1_sub_fp_4_10 <= 1 << index_trunc_4_10;
        l1_valid_4_10 <= 1;
    end
    l1_sub_fp_4_11 <= 0;
    l1_valid_4_11 <= 0;
    if(din_valid_4_11)begin
        l1_sub_fp_4_11 <= 1 << index_trunc_4_11;
        l1_valid_4_11 <= 1;
    end
    l1_sub_fp_4_12 <= 0;
    l1_valid_4_12 <= 0;
    if(din_valid_4_12)begin
        l1_sub_fp_4_12 <= 1 << index_trunc_4_12;
        l1_valid_4_12 <= 1;
    end
    l1_sub_fp_4_13 <= 0;
    l1_valid_4_13 <= 0;
    if(din_valid_4_13)begin
        l1_sub_fp_4_13 <= 1 << index_trunc_4_13;
        l1_valid_4_13 <= 1;
    end
    l1_sub_fp_4_14 <= 0;
    l1_valid_4_14 <= 0;
    if(din_valid_4_14)begin
        l1_sub_fp_4_14 <= 1 << index_trunc_4_14;
        l1_valid_4_14 <= 1;
    end
    l1_sub_fp_4_15 <= 0;
    l1_valid_4_15 <= 0;
    if(din_valid_4_15)begin
        l1_sub_fp_4_15 <= 1 << index_trunc_4_15;
        l1_valid_4_15 <= 1;
    end
    l1_sub_fp_5_0 <= 0;
    l1_valid_5_0 <= 0;
    if(din_valid_5_0)begin
        l1_sub_fp_5_0 <= 1 << index_trunc_5_0;
        l1_valid_5_0 <= 1;
    end
    l1_sub_fp_5_1 <= 0;
    l1_valid_5_1 <= 0;
    if(din_valid_5_1)begin
        l1_sub_fp_5_1 <= 1 << index_trunc_5_1;
        l1_valid_5_1 <= 1;
    end
    l1_sub_fp_5_2 <= 0;
    l1_valid_5_2 <= 0;
    if(din_valid_5_2)begin
        l1_sub_fp_5_2 <= 1 << index_trunc_5_2;
        l1_valid_5_2 <= 1;
    end
    l1_sub_fp_5_3 <= 0;
    l1_valid_5_3 <= 0;
    if(din_valid_5_3)begin
        l1_sub_fp_5_3 <= 1 << index_trunc_5_3;
        l1_valid_5_3 <= 1;
    end
    l1_sub_fp_5_4 <= 0;
    l1_valid_5_4 <= 0;
    if(din_valid_5_4)begin
        l1_sub_fp_5_4 <= 1 << index_trunc_5_4;
        l1_valid_5_4 <= 1;
    end
    l1_sub_fp_5_5 <= 0;
    l1_valid_5_5 <= 0;
    if(din_valid_5_5)begin
        l1_sub_fp_5_5 <= 1 << index_trunc_5_5;
        l1_valid_5_5 <= 1;
    end
    l1_sub_fp_5_6 <= 0;
    l1_valid_5_6 <= 0;
    if(din_valid_5_6)begin
        l1_sub_fp_5_6 <= 1 << index_trunc_5_6;
        l1_valid_5_6 <= 1;
    end
    l1_sub_fp_5_7 <= 0;
    l1_valid_5_7 <= 0;
    if(din_valid_5_7)begin
        l1_sub_fp_5_7 <= 1 << index_trunc_5_7;
        l1_valid_5_7 <= 1;
    end
    l1_sub_fp_5_8 <= 0;
    l1_valid_5_8 <= 0;
    if(din_valid_5_8)begin
        l1_sub_fp_5_8 <= 1 << index_trunc_5_8;
        l1_valid_5_8 <= 1;
    end
    l1_sub_fp_5_9 <= 0;
    l1_valid_5_9 <= 0;
    if(din_valid_5_9)begin
        l1_sub_fp_5_9 <= 1 << index_trunc_5_9;
        l1_valid_5_9 <= 1;
    end
    l1_sub_fp_5_10 <= 0;
    l1_valid_5_10 <= 0;
    if(din_valid_5_10)begin
        l1_sub_fp_5_10 <= 1 << index_trunc_5_10;
        l1_valid_5_10 <= 1;
    end
    l1_sub_fp_5_11 <= 0;
    l1_valid_5_11 <= 0;
    if(din_valid_5_11)begin
        l1_sub_fp_5_11 <= 1 << index_trunc_5_11;
        l1_valid_5_11 <= 1;
    end
    l1_sub_fp_5_12 <= 0;
    l1_valid_5_12 <= 0;
    if(din_valid_5_12)begin
        l1_sub_fp_5_12 <= 1 << index_trunc_5_12;
        l1_valid_5_12 <= 1;
    end
    l1_sub_fp_5_13 <= 0;
    l1_valid_5_13 <= 0;
    if(din_valid_5_13)begin
        l1_sub_fp_5_13 <= 1 << index_trunc_5_13;
        l1_valid_5_13 <= 1;
    end
    l1_sub_fp_5_14 <= 0;
    l1_valid_5_14 <= 0;
    if(din_valid_5_14)begin
        l1_sub_fp_5_14 <= 1 << index_trunc_5_14;
        l1_valid_5_14 <= 1;
    end
    l1_sub_fp_5_15 <= 0;
    l1_valid_5_15 <= 0;
    if(din_valid_5_15)begin
        l1_sub_fp_5_15 <= 1 << index_trunc_5_15;
        l1_valid_5_15 <= 1;
    end
    l1_sub_fp_6_0 <= 0;
    l1_valid_6_0 <= 0;
    if(din_valid_6_0)begin
        l1_sub_fp_6_0 <= 1 << index_trunc_6_0;
        l1_valid_6_0 <= 1;
    end
    l1_sub_fp_6_1 <= 0;
    l1_valid_6_1 <= 0;
    if(din_valid_6_1)begin
        l1_sub_fp_6_1 <= 1 << index_trunc_6_1;
        l1_valid_6_1 <= 1;
    end
    l1_sub_fp_6_2 <= 0;
    l1_valid_6_2 <= 0;
    if(din_valid_6_2)begin
        l1_sub_fp_6_2 <= 1 << index_trunc_6_2;
        l1_valid_6_2 <= 1;
    end
    l1_sub_fp_6_3 <= 0;
    l1_valid_6_3 <= 0;
    if(din_valid_6_3)begin
        l1_sub_fp_6_3 <= 1 << index_trunc_6_3;
        l1_valid_6_3 <= 1;
    end
    l1_sub_fp_6_4 <= 0;
    l1_valid_6_4 <= 0;
    if(din_valid_6_4)begin
        l1_sub_fp_6_4 <= 1 << index_trunc_6_4;
        l1_valid_6_4 <= 1;
    end
    l1_sub_fp_6_5 <= 0;
    l1_valid_6_5 <= 0;
    if(din_valid_6_5)begin
        l1_sub_fp_6_5 <= 1 << index_trunc_6_5;
        l1_valid_6_5 <= 1;
    end
    l1_sub_fp_6_6 <= 0;
    l1_valid_6_6 <= 0;
    if(din_valid_6_6)begin
        l1_sub_fp_6_6 <= 1 << index_trunc_6_6;
        l1_valid_6_6 <= 1;
    end
    l1_sub_fp_6_7 <= 0;
    l1_valid_6_7 <= 0;
    if(din_valid_6_7)begin
        l1_sub_fp_6_7 <= 1 << index_trunc_6_7;
        l1_valid_6_7 <= 1;
    end
    l1_sub_fp_6_8 <= 0;
    l1_valid_6_8 <= 0;
    if(din_valid_6_8)begin
        l1_sub_fp_6_8 <= 1 << index_trunc_6_8;
        l1_valid_6_8 <= 1;
    end
    l1_sub_fp_6_9 <= 0;
    l1_valid_6_9 <= 0;
    if(din_valid_6_9)begin
        l1_sub_fp_6_9 <= 1 << index_trunc_6_9;
        l1_valid_6_9 <= 1;
    end
    l1_sub_fp_6_10 <= 0;
    l1_valid_6_10 <= 0;
    if(din_valid_6_10)begin
        l1_sub_fp_6_10 <= 1 << index_trunc_6_10;
        l1_valid_6_10 <= 1;
    end
    l1_sub_fp_6_11 <= 0;
    l1_valid_6_11 <= 0;
    if(din_valid_6_11)begin
        l1_sub_fp_6_11 <= 1 << index_trunc_6_11;
        l1_valid_6_11 <= 1;
    end
    l1_sub_fp_6_12 <= 0;
    l1_valid_6_12 <= 0;
    if(din_valid_6_12)begin
        l1_sub_fp_6_12 <= 1 << index_trunc_6_12;
        l1_valid_6_12 <= 1;
    end
    l1_sub_fp_6_13 <= 0;
    l1_valid_6_13 <= 0;
    if(din_valid_6_13)begin
        l1_sub_fp_6_13 <= 1 << index_trunc_6_13;
        l1_valid_6_13 <= 1;
    end
    l1_sub_fp_6_14 <= 0;
    l1_valid_6_14 <= 0;
    if(din_valid_6_14)begin
        l1_sub_fp_6_14 <= 1 << index_trunc_6_14;
        l1_valid_6_14 <= 1;
    end
    l1_sub_fp_6_15 <= 0;
    l1_valid_6_15 <= 0;
    if(din_valid_6_15)begin
        l1_sub_fp_6_15 <= 1 << index_trunc_6_15;
        l1_valid_6_15 <= 1;
    end
    l1_sub_fp_7_0 <= 0;
    l1_valid_7_0 <= 0;
    if(din_valid_7_0)begin
        l1_sub_fp_7_0 <= 1 << index_trunc_7_0;
        l1_valid_7_0 <= 1;
    end
    l1_sub_fp_7_1 <= 0;
    l1_valid_7_1 <= 0;
    if(din_valid_7_1)begin
        l1_sub_fp_7_1 <= 1 << index_trunc_7_1;
        l1_valid_7_1 <= 1;
    end
    l1_sub_fp_7_2 <= 0;
    l1_valid_7_2 <= 0;
    if(din_valid_7_2)begin
        l1_sub_fp_7_2 <= 1 << index_trunc_7_2;
        l1_valid_7_2 <= 1;
    end
    l1_sub_fp_7_3 <= 0;
    l1_valid_7_3 <= 0;
    if(din_valid_7_3)begin
        l1_sub_fp_7_3 <= 1 << index_trunc_7_3;
        l1_valid_7_3 <= 1;
    end
    l1_sub_fp_7_4 <= 0;
    l1_valid_7_4 <= 0;
    if(din_valid_7_4)begin
        l1_sub_fp_7_4 <= 1 << index_trunc_7_4;
        l1_valid_7_4 <= 1;
    end
    l1_sub_fp_7_5 <= 0;
    l1_valid_7_5 <= 0;
    if(din_valid_7_5)begin
        l1_sub_fp_7_5 <= 1 << index_trunc_7_5;
        l1_valid_7_5 <= 1;
    end
    l1_sub_fp_7_6 <= 0;
    l1_valid_7_6 <= 0;
    if(din_valid_7_6)begin
        l1_sub_fp_7_6 <= 1 << index_trunc_7_6;
        l1_valid_7_6 <= 1;
    end
    l1_sub_fp_7_7 <= 0;
    l1_valid_7_7 <= 0;
    if(din_valid_7_7)begin
        l1_sub_fp_7_7 <= 1 << index_trunc_7_7;
        l1_valid_7_7 <= 1;
    end
    l1_sub_fp_7_8 <= 0;
    l1_valid_7_8 <= 0;
    if(din_valid_7_8)begin
        l1_sub_fp_7_8 <= 1 << index_trunc_7_8;
        l1_valid_7_8 <= 1;
    end
    l1_sub_fp_7_9 <= 0;
    l1_valid_7_9 <= 0;
    if(din_valid_7_9)begin
        l1_sub_fp_7_9 <= 1 << index_trunc_7_9;
        l1_valid_7_9 <= 1;
    end
    l1_sub_fp_7_10 <= 0;
    l1_valid_7_10 <= 0;
    if(din_valid_7_10)begin
        l1_sub_fp_7_10 <= 1 << index_trunc_7_10;
        l1_valid_7_10 <= 1;
    end
    l1_sub_fp_7_11 <= 0;
    l1_valid_7_11 <= 0;
    if(din_valid_7_11)begin
        l1_sub_fp_7_11 <= 1 << index_trunc_7_11;
        l1_valid_7_11 <= 1;
    end
    l1_sub_fp_7_12 <= 0;
    l1_valid_7_12 <= 0;
    if(din_valid_7_12)begin
        l1_sub_fp_7_12 <= 1 << index_trunc_7_12;
        l1_valid_7_12 <= 1;
    end
    l1_sub_fp_7_13 <= 0;
    l1_valid_7_13 <= 0;
    if(din_valid_7_13)begin
        l1_sub_fp_7_13 <= 1 << index_trunc_7_13;
        l1_valid_7_13 <= 1;
    end
    l1_sub_fp_7_14 <= 0;
    l1_valid_7_14 <= 0;
    if(din_valid_7_14)begin
        l1_sub_fp_7_14 <= 1 << index_trunc_7_14;
        l1_valid_7_14 <= 1;
    end
    l1_sub_fp_7_15 <= 0;
    l1_valid_7_15 <= 0;
    if(din_valid_7_15)begin
        l1_sub_fp_7_15 <= 1 << index_trunc_7_15;
        l1_valid_7_15 <= 1;
    end
end

//Layer 2
always@(posedge clk)begin
    l2_sub_fp_0_0 <= 0;
    l2_valid_0_0  <= 0;
    if(l1_valid_0_0 | l1_valid_0_1)begin
        l2_sub_fp_0_0 <= l1_sub_fp_0_0 | l1_sub_fp_0_1;
        l2_valid_0_0 <= 1;
    end
    l2_sub_fp_0_1 <= 0;
    l2_valid_0_1  <= 0;
    if(l1_valid_0_2 | l1_valid_0_3)begin
        l2_sub_fp_0_1 <= l1_sub_fp_0_2 | l1_sub_fp_0_3;
        l2_valid_0_1 <= 1;
    end
    l2_sub_fp_0_2 <= 0;
    l2_valid_0_2  <= 0;
    if(l1_valid_0_4 | l1_valid_0_5)begin
        l2_sub_fp_0_2 <= l1_sub_fp_0_4 | l1_sub_fp_0_5;
        l2_valid_0_2 <= 1;
    end
    l2_sub_fp_0_3 <= 0;
    l2_valid_0_3  <= 0;
    if(l1_valid_0_6 | l1_valid_0_7)begin
        l2_sub_fp_0_3 <= l1_sub_fp_0_6 | l1_sub_fp_0_7;
        l2_valid_0_3 <= 1;
    end
    l2_sub_fp_0_4 <= 0;
    l2_valid_0_4  <= 0;
    if(l1_valid_0_8 | l1_valid_0_9)begin
        l2_sub_fp_0_4 <= l1_sub_fp_0_8 | l1_sub_fp_0_9;
        l2_valid_0_4 <= 1;
    end
    l2_sub_fp_0_5 <= 0;
    l2_valid_0_5  <= 0;
    if(l1_valid_0_10 | l1_valid_0_11)begin
        l2_sub_fp_0_5 <= l1_sub_fp_0_10 | l1_sub_fp_0_11;
        l2_valid_0_5 <= 1;
    end
    l2_sub_fp_0_6 <= 0;
    l2_valid_0_6  <= 0;
    if(l1_valid_0_12 | l1_valid_0_13)begin
        l2_sub_fp_0_6 <= l1_sub_fp_0_12 | l1_sub_fp_0_13;
        l2_valid_0_6 <= 1;
    end
    l2_sub_fp_0_7 <= 0;
    l2_valid_0_7  <= 0;
    if(l1_valid_0_14 | l1_valid_0_15)begin
        l2_sub_fp_0_7 <= l1_sub_fp_0_14 | l1_sub_fp_0_15;
        l2_valid_0_7 <= 1;
    end
    l2_sub_fp_1_0 <= 0;
    l2_valid_1_0  <= 0;
    if(l1_valid_1_0 | l1_valid_1_1)begin
        l2_sub_fp_1_0 <= l1_sub_fp_1_0 | l1_sub_fp_1_1;
        l2_valid_1_0 <= 1;
    end
    l2_sub_fp_1_1 <= 0;
    l2_valid_1_1  <= 0;
    if(l1_valid_1_2 | l1_valid_1_3)begin
        l2_sub_fp_1_1 <= l1_sub_fp_1_2 | l1_sub_fp_1_3;
        l2_valid_1_1 <= 1;
    end
    l2_sub_fp_1_2 <= 0;
    l2_valid_1_2  <= 0;
    if(l1_valid_1_4 | l1_valid_1_5)begin
        l2_sub_fp_1_2 <= l1_sub_fp_1_4 | l1_sub_fp_1_5;
        l2_valid_1_2 <= 1;
    end
    l2_sub_fp_1_3 <= 0;
    l2_valid_1_3  <= 0;
    if(l1_valid_1_6 | l1_valid_1_7)begin
        l2_sub_fp_1_3 <= l1_sub_fp_1_6 | l1_sub_fp_1_7;
        l2_valid_1_3 <= 1;
    end
    l2_sub_fp_1_4 <= 0;
    l2_valid_1_4  <= 0;
    if(l1_valid_1_8 | l1_valid_1_9)begin
        l2_sub_fp_1_4 <= l1_sub_fp_1_8 | l1_sub_fp_1_9;
        l2_valid_1_4 <= 1;
    end
    l2_sub_fp_1_5 <= 0;
    l2_valid_1_5  <= 0;
    if(l1_valid_1_10 | l1_valid_1_11)begin
        l2_sub_fp_1_5 <= l1_sub_fp_1_10 | l1_sub_fp_1_11;
        l2_valid_1_5 <= 1;
    end
    l2_sub_fp_1_6 <= 0;
    l2_valid_1_6  <= 0;
    if(l1_valid_1_12 | l1_valid_1_13)begin
        l2_sub_fp_1_6 <= l1_sub_fp_1_12 | l1_sub_fp_1_13;
        l2_valid_1_6 <= 1;
    end
    l2_sub_fp_1_7 <= 0;
    l2_valid_1_7  <= 0;
    if(l1_valid_1_14 | l1_valid_1_15)begin
        l2_sub_fp_1_7 <= l1_sub_fp_1_14 | l1_sub_fp_1_15;
        l2_valid_1_7 <= 1;
    end
    l2_sub_fp_2_0 <= 0;
    l2_valid_2_0  <= 0;
    if(l1_valid_2_0 | l1_valid_2_1)begin
        l2_sub_fp_2_0 <= l1_sub_fp_2_0 | l1_sub_fp_2_1;
        l2_valid_2_0 <= 1;
    end
    l2_sub_fp_2_1 <= 0;
    l2_valid_2_1  <= 0;
    if(l1_valid_2_2 | l1_valid_2_3)begin
        l2_sub_fp_2_1 <= l1_sub_fp_2_2 | l1_sub_fp_2_3;
        l2_valid_2_1 <= 1;
    end
    l2_sub_fp_2_2 <= 0;
    l2_valid_2_2  <= 0;
    if(l1_valid_2_4 | l1_valid_2_5)begin
        l2_sub_fp_2_2 <= l1_sub_fp_2_4 | l1_sub_fp_2_5;
        l2_valid_2_2 <= 1;
    end
    l2_sub_fp_2_3 <= 0;
    l2_valid_2_3  <= 0;
    if(l1_valid_2_6 | l1_valid_2_7)begin
        l2_sub_fp_2_3 <= l1_sub_fp_2_6 | l1_sub_fp_2_7;
        l2_valid_2_3 <= 1;
    end
    l2_sub_fp_2_4 <= 0;
    l2_valid_2_4  <= 0;
    if(l1_valid_2_8 | l1_valid_2_9)begin
        l2_sub_fp_2_4 <= l1_sub_fp_2_8 | l1_sub_fp_2_9;
        l2_valid_2_4 <= 1;
    end
    l2_sub_fp_2_5 <= 0;
    l2_valid_2_5  <= 0;
    if(l1_valid_2_10 | l1_valid_2_11)begin
        l2_sub_fp_2_5 <= l1_sub_fp_2_10 | l1_sub_fp_2_11;
        l2_valid_2_5 <= 1;
    end
    l2_sub_fp_2_6 <= 0;
    l2_valid_2_6  <= 0;
    if(l1_valid_2_12 | l1_valid_2_13)begin
        l2_sub_fp_2_6 <= l1_sub_fp_2_12 | l1_sub_fp_2_13;
        l2_valid_2_6 <= 1;
    end
    l2_sub_fp_2_7 <= 0;
    l2_valid_2_7  <= 0;
    if(l1_valid_2_14 | l1_valid_2_15)begin
        l2_sub_fp_2_7 <= l1_sub_fp_2_14 | l1_sub_fp_2_15;
        l2_valid_2_7 <= 1;
    end
    l2_sub_fp_3_0 <= 0;
    l2_valid_3_0  <= 0;
    if(l1_valid_3_0 | l1_valid_3_1)begin
        l2_sub_fp_3_0 <= l1_sub_fp_3_0 | l1_sub_fp_3_1;
        l2_valid_3_0 <= 1;
    end
    l2_sub_fp_3_1 <= 0;
    l2_valid_3_1  <= 0;
    if(l1_valid_3_2 | l1_valid_3_3)begin
        l2_sub_fp_3_1 <= l1_sub_fp_3_2 | l1_sub_fp_3_3;
        l2_valid_3_1 <= 1;
    end
    l2_sub_fp_3_2 <= 0;
    l2_valid_3_2  <= 0;
    if(l1_valid_3_4 | l1_valid_3_5)begin
        l2_sub_fp_3_2 <= l1_sub_fp_3_4 | l1_sub_fp_3_5;
        l2_valid_3_2 <= 1;
    end
    l2_sub_fp_3_3 <= 0;
    l2_valid_3_3  <= 0;
    if(l1_valid_3_6 | l1_valid_3_7)begin
        l2_sub_fp_3_3 <= l1_sub_fp_3_6 | l1_sub_fp_3_7;
        l2_valid_3_3 <= 1;
    end
    l2_sub_fp_3_4 <= 0;
    l2_valid_3_4  <= 0;
    if(l1_valid_3_8 | l1_valid_3_9)begin
        l2_sub_fp_3_4 <= l1_sub_fp_3_8 | l1_sub_fp_3_9;
        l2_valid_3_4 <= 1;
    end
    l2_sub_fp_3_5 <= 0;
    l2_valid_3_5  <= 0;
    if(l1_valid_3_10 | l1_valid_3_11)begin
        l2_sub_fp_3_5 <= l1_sub_fp_3_10 | l1_sub_fp_3_11;
        l2_valid_3_5 <= 1;
    end
    l2_sub_fp_3_6 <= 0;
    l2_valid_3_6  <= 0;
    if(l1_valid_3_12 | l1_valid_3_13)begin
        l2_sub_fp_3_6 <= l1_sub_fp_3_12 | l1_sub_fp_3_13;
        l2_valid_3_6 <= 1;
    end
    l2_sub_fp_3_7 <= 0;
    l2_valid_3_7  <= 0;
    if(l1_valid_3_14 | l1_valid_3_15)begin
        l2_sub_fp_3_7 <= l1_sub_fp_3_14 | l1_sub_fp_3_15;
        l2_valid_3_7 <= 1;
    end
    l2_sub_fp_4_0 <= 0;
    l2_valid_4_0  <= 0;
    if(l1_valid_4_0 | l1_valid_4_1)begin
        l2_sub_fp_4_0 <= l1_sub_fp_4_0 | l1_sub_fp_4_1;
        l2_valid_4_0 <= 1;
    end
    l2_sub_fp_4_1 <= 0;
    l2_valid_4_1  <= 0;
    if(l1_valid_4_2 | l1_valid_4_3)begin
        l2_sub_fp_4_1 <= l1_sub_fp_4_2 | l1_sub_fp_4_3;
        l2_valid_4_1 <= 1;
    end
    l2_sub_fp_4_2 <= 0;
    l2_valid_4_2  <= 0;
    if(l1_valid_4_4 | l1_valid_4_5)begin
        l2_sub_fp_4_2 <= l1_sub_fp_4_4 | l1_sub_fp_4_5;
        l2_valid_4_2 <= 1;
    end
    l2_sub_fp_4_3 <= 0;
    l2_valid_4_3  <= 0;
    if(l1_valid_4_6 | l1_valid_4_7)begin
        l2_sub_fp_4_3 <= l1_sub_fp_4_6 | l1_sub_fp_4_7;
        l2_valid_4_3 <= 1;
    end
    l2_sub_fp_4_4 <= 0;
    l2_valid_4_4  <= 0;
    if(l1_valid_4_8 | l1_valid_4_9)begin
        l2_sub_fp_4_4 <= l1_sub_fp_4_8 | l1_sub_fp_4_9;
        l2_valid_4_4 <= 1;
    end
    l2_sub_fp_4_5 <= 0;
    l2_valid_4_5  <= 0;
    if(l1_valid_4_10 | l1_valid_4_11)begin
        l2_sub_fp_4_5 <= l1_sub_fp_4_10 | l1_sub_fp_4_11;
        l2_valid_4_5 <= 1;
    end
    l2_sub_fp_4_6 <= 0;
    l2_valid_4_6  <= 0;
    if(l1_valid_4_12 | l1_valid_4_13)begin
        l2_sub_fp_4_6 <= l1_sub_fp_4_12 | l1_sub_fp_4_13;
        l2_valid_4_6 <= 1;
    end
    l2_sub_fp_4_7 <= 0;
    l2_valid_4_7  <= 0;
    if(l1_valid_4_14 | l1_valid_4_15)begin
        l2_sub_fp_4_7 <= l1_sub_fp_4_14 | l1_sub_fp_4_15;
        l2_valid_4_7 <= 1;
    end
    l2_sub_fp_5_0 <= 0;
    l2_valid_5_0  <= 0;
    if(l1_valid_5_0 | l1_valid_5_1)begin
        l2_sub_fp_5_0 <= l1_sub_fp_5_0 | l1_sub_fp_5_1;
        l2_valid_5_0 <= 1;
    end
    l2_sub_fp_5_1 <= 0;
    l2_valid_5_1  <= 0;
    if(l1_valid_5_2 | l1_valid_5_3)begin
        l2_sub_fp_5_1 <= l1_sub_fp_5_2 | l1_sub_fp_5_3;
        l2_valid_5_1 <= 1;
    end
    l2_sub_fp_5_2 <= 0;
    l2_valid_5_2  <= 0;
    if(l1_valid_5_4 | l1_valid_5_5)begin
        l2_sub_fp_5_2 <= l1_sub_fp_5_4 | l1_sub_fp_5_5;
        l2_valid_5_2 <= 1;
    end
    l2_sub_fp_5_3 <= 0;
    l2_valid_5_3  <= 0;
    if(l1_valid_5_6 | l1_valid_5_7)begin
        l2_sub_fp_5_3 <= l1_sub_fp_5_6 | l1_sub_fp_5_7;
        l2_valid_5_3 <= 1;
    end
    l2_sub_fp_5_4 <= 0;
    l2_valid_5_4  <= 0;
    if(l1_valid_5_8 | l1_valid_5_9)begin
        l2_sub_fp_5_4 <= l1_sub_fp_5_8 | l1_sub_fp_5_9;
        l2_valid_5_4 <= 1;
    end
    l2_sub_fp_5_5 <= 0;
    l2_valid_5_5  <= 0;
    if(l1_valid_5_10 | l1_valid_5_11)begin
        l2_sub_fp_5_5 <= l1_sub_fp_5_10 | l1_sub_fp_5_11;
        l2_valid_5_5 <= 1;
    end
    l2_sub_fp_5_6 <= 0;
    l2_valid_5_6  <= 0;
    if(l1_valid_5_12 | l1_valid_5_13)begin
        l2_sub_fp_5_6 <= l1_sub_fp_5_12 | l1_sub_fp_5_13;
        l2_valid_5_6 <= 1;
    end
    l2_sub_fp_5_7 <= 0;
    l2_valid_5_7  <= 0;
    if(l1_valid_5_14 | l1_valid_5_15)begin
        l2_sub_fp_5_7 <= l1_sub_fp_5_14 | l1_sub_fp_5_15;
        l2_valid_5_7 <= 1;
    end
    l2_sub_fp_6_0 <= 0;
    l2_valid_6_0  <= 0;
    if(l1_valid_6_0 | l1_valid_6_1)begin
        l2_sub_fp_6_0 <= l1_sub_fp_6_0 | l1_sub_fp_6_1;
        l2_valid_6_0 <= 1;
    end
    l2_sub_fp_6_1 <= 0;
    l2_valid_6_1  <= 0;
    if(l1_valid_6_2 | l1_valid_6_3)begin
        l2_sub_fp_6_1 <= l1_sub_fp_6_2 | l1_sub_fp_6_3;
        l2_valid_6_1 <= 1;
    end
    l2_sub_fp_6_2 <= 0;
    l2_valid_6_2  <= 0;
    if(l1_valid_6_4 | l1_valid_6_5)begin
        l2_sub_fp_6_2 <= l1_sub_fp_6_4 | l1_sub_fp_6_5;
        l2_valid_6_2 <= 1;
    end
    l2_sub_fp_6_3 <= 0;
    l2_valid_6_3  <= 0;
    if(l1_valid_6_6 | l1_valid_6_7)begin
        l2_sub_fp_6_3 <= l1_sub_fp_6_6 | l1_sub_fp_6_7;
        l2_valid_6_3 <= 1;
    end
    l2_sub_fp_6_4 <= 0;
    l2_valid_6_4  <= 0;
    if(l1_valid_6_8 | l1_valid_6_9)begin
        l2_sub_fp_6_4 <= l1_sub_fp_6_8 | l1_sub_fp_6_9;
        l2_valid_6_4 <= 1;
    end
    l2_sub_fp_6_5 <= 0;
    l2_valid_6_5  <= 0;
    if(l1_valid_6_10 | l1_valid_6_11)begin
        l2_sub_fp_6_5 <= l1_sub_fp_6_10 | l1_sub_fp_6_11;
        l2_valid_6_5 <= 1;
    end
    l2_sub_fp_6_6 <= 0;
    l2_valid_6_6  <= 0;
    if(l1_valid_6_12 | l1_valid_6_13)begin
        l2_sub_fp_6_6 <= l1_sub_fp_6_12 | l1_sub_fp_6_13;
        l2_valid_6_6 <= 1;
    end
    l2_sub_fp_6_7 <= 0;
    l2_valid_6_7  <= 0;
    if(l1_valid_6_14 | l1_valid_6_15)begin
        l2_sub_fp_6_7 <= l1_sub_fp_6_14 | l1_sub_fp_6_15;
        l2_valid_6_7 <= 1;
    end
    l2_sub_fp_7_0 <= 0;
    l2_valid_7_0  <= 0;
    if(l1_valid_7_0 | l1_valid_7_1)begin
        l2_sub_fp_7_0 <= l1_sub_fp_7_0 | l1_sub_fp_7_1;
        l2_valid_7_0 <= 1;
    end
    l2_sub_fp_7_1 <= 0;
    l2_valid_7_1  <= 0;
    if(l1_valid_7_2 | l1_valid_7_3)begin
        l2_sub_fp_7_1 <= l1_sub_fp_7_2 | l1_sub_fp_7_3;
        l2_valid_7_1 <= 1;
    end
    l2_sub_fp_7_2 <= 0;
    l2_valid_7_2  <= 0;
    if(l1_valid_7_4 | l1_valid_7_5)begin
        l2_sub_fp_7_2 <= l1_sub_fp_7_4 | l1_sub_fp_7_5;
        l2_valid_7_2 <= 1;
    end
    l2_sub_fp_7_3 <= 0;
    l2_valid_7_3  <= 0;
    if(l1_valid_7_6 | l1_valid_7_7)begin
        l2_sub_fp_7_3 <= l1_sub_fp_7_6 | l1_sub_fp_7_7;
        l2_valid_7_3 <= 1;
    end
    l2_sub_fp_7_4 <= 0;
    l2_valid_7_4  <= 0;
    if(l1_valid_7_8 | l1_valid_7_9)begin
        l2_sub_fp_7_4 <= l1_sub_fp_7_8 | l1_sub_fp_7_9;
        l2_valid_7_4 <= 1;
    end
    l2_sub_fp_7_5 <= 0;
    l2_valid_7_5  <= 0;
    if(l1_valid_7_10 | l1_valid_7_11)begin
        l2_sub_fp_7_5 <= l1_sub_fp_7_10 | l1_sub_fp_7_11;
        l2_valid_7_5 <= 1;
    end
    l2_sub_fp_7_6 <= 0;
    l2_valid_7_6  <= 0;
    if(l1_valid_7_12 | l1_valid_7_13)begin
        l2_sub_fp_7_6 <= l1_sub_fp_7_12 | l1_sub_fp_7_13;
        l2_valid_7_6 <= 1;
    end
    l2_sub_fp_7_7 <= 0;
    l2_valid_7_7  <= 0;
    if(l1_valid_7_14 | l1_valid_7_15)begin
        l2_sub_fp_7_7 <= l1_sub_fp_7_14 | l1_sub_fp_7_15;
        l2_valid_7_7 <= 1;
    end
end

//Layer 3
always@(posedge clk)begin
    l3_sub_fp_0_0 <= 0;
    l3_valid_0_0  <= 0;
    if(l2_valid_0_0 | l2_valid_0_1)begin
        l3_sub_fp_0_0 <= l2_sub_fp_0_0 | l2_sub_fp_0_1;
        l3_valid_0_0 <= 1;
    end
    l3_sub_fp_0_1 <= 0;
    l3_valid_0_1  <= 0;
    if(l2_valid_0_2 | l2_valid_0_3)begin
        l3_sub_fp_0_1 <= l2_sub_fp_0_2 | l2_sub_fp_0_3;
        l3_valid_0_1 <= 1;
    end
    l3_sub_fp_0_2 <= 0;
    l3_valid_0_2  <= 0;
    if(l2_valid_0_4 | l2_valid_0_5)begin
        l3_sub_fp_0_2 <= l2_sub_fp_0_4 | l2_sub_fp_0_5;
        l3_valid_0_2 <= 1;
    end
    l3_sub_fp_0_3 <= 0;
    l3_valid_0_3  <= 0;
    if(l2_valid_0_6 | l2_valid_0_7)begin
        l3_sub_fp_0_3 <= l2_sub_fp_0_6 | l2_sub_fp_0_7;
        l3_valid_0_3 <= 1;
    end
    l3_sub_fp_1_0 <= 0;
    l3_valid_1_0  <= 0;
    if(l2_valid_1_0 | l2_valid_1_1)begin
        l3_sub_fp_1_0 <= l2_sub_fp_1_0 | l2_sub_fp_1_1;
        l3_valid_1_0 <= 1;
    end
    l3_sub_fp_1_1 <= 0;
    l3_valid_1_1  <= 0;
    if(l2_valid_1_2 | l2_valid_1_3)begin
        l3_sub_fp_1_1 <= l2_sub_fp_1_2 | l2_sub_fp_1_3;
        l3_valid_1_1 <= 1;
    end
    l3_sub_fp_1_2 <= 0;
    l3_valid_1_2  <= 0;
    if(l2_valid_1_4 | l2_valid_1_5)begin
        l3_sub_fp_1_2 <= l2_sub_fp_1_4 | l2_sub_fp_1_5;
        l3_valid_1_2 <= 1;
    end
    l3_sub_fp_1_3 <= 0;
    l3_valid_1_3  <= 0;
    if(l2_valid_1_6 | l2_valid_1_7)begin
        l3_sub_fp_1_3 <= l2_sub_fp_1_6 | l2_sub_fp_1_7;
        l3_valid_1_3 <= 1;
    end
    l3_sub_fp_2_0 <= 0;
    l3_valid_2_0  <= 0;
    if(l2_valid_2_0 | l2_valid_2_1)begin
        l3_sub_fp_2_0 <= l2_sub_fp_2_0 | l2_sub_fp_2_1;
        l3_valid_2_0 <= 1;
    end
    l3_sub_fp_2_1 <= 0;
    l3_valid_2_1  <= 0;
    if(l2_valid_2_2 | l2_valid_2_3)begin
        l3_sub_fp_2_1 <= l2_sub_fp_2_2 | l2_sub_fp_2_3;
        l3_valid_2_1 <= 1;
    end
    l3_sub_fp_2_2 <= 0;
    l3_valid_2_2  <= 0;
    if(l2_valid_2_4 | l2_valid_2_5)begin
        l3_sub_fp_2_2 <= l2_sub_fp_2_4 | l2_sub_fp_2_5;
        l3_valid_2_2 <= 1;
    end
    l3_sub_fp_2_3 <= 0;
    l3_valid_2_3  <= 0;
    if(l2_valid_2_6 | l2_valid_2_7)begin
        l3_sub_fp_2_3 <= l2_sub_fp_2_6 | l2_sub_fp_2_7;
        l3_valid_2_3 <= 1;
    end
    l3_sub_fp_3_0 <= 0;
    l3_valid_3_0  <= 0;
    if(l2_valid_3_0 | l2_valid_3_1)begin
        l3_sub_fp_3_0 <= l2_sub_fp_3_0 | l2_sub_fp_3_1;
        l3_valid_3_0 <= 1;
    end
    l3_sub_fp_3_1 <= 0;
    l3_valid_3_1  <= 0;
    if(l2_valid_3_2 | l2_valid_3_3)begin
        l3_sub_fp_3_1 <= l2_sub_fp_3_2 | l2_sub_fp_3_3;
        l3_valid_3_1 <= 1;
    end
    l3_sub_fp_3_2 <= 0;
    l3_valid_3_2  <= 0;
    if(l2_valid_3_4 | l2_valid_3_5)begin
        l3_sub_fp_3_2 <= l2_sub_fp_3_4 | l2_sub_fp_3_5;
        l3_valid_3_2 <= 1;
    end
    l3_sub_fp_3_3 <= 0;
    l3_valid_3_3  <= 0;
    if(l2_valid_3_6 | l2_valid_3_7)begin
        l3_sub_fp_3_3 <= l2_sub_fp_3_6 | l2_sub_fp_3_7;
        l3_valid_3_3 <= 1;
    end
    l3_sub_fp_4_0 <= 0;
    l3_valid_4_0  <= 0;
    if(l2_valid_4_0 | l2_valid_4_1)begin
        l3_sub_fp_4_0 <= l2_sub_fp_4_0 | l2_sub_fp_4_1;
        l3_valid_4_0 <= 1;
    end
    l3_sub_fp_4_1 <= 0;
    l3_valid_4_1  <= 0;
    if(l2_valid_4_2 | l2_valid_4_3)begin
        l3_sub_fp_4_1 <= l2_sub_fp_4_2 | l2_sub_fp_4_3;
        l3_valid_4_1 <= 1;
    end
    l3_sub_fp_4_2 <= 0;
    l3_valid_4_2  <= 0;
    if(l2_valid_4_4 | l2_valid_4_5)begin
        l3_sub_fp_4_2 <= l2_sub_fp_4_4 | l2_sub_fp_4_5;
        l3_valid_4_2 <= 1;
    end
    l3_sub_fp_4_3 <= 0;
    l3_valid_4_3  <= 0;
    if(l2_valid_4_6 | l2_valid_4_7)begin
        l3_sub_fp_4_3 <= l2_sub_fp_4_6 | l2_sub_fp_4_7;
        l3_valid_4_3 <= 1;
    end
    l3_sub_fp_5_0 <= 0;
    l3_valid_5_0  <= 0;
    if(l2_valid_5_0 | l2_valid_5_1)begin
        l3_sub_fp_5_0 <= l2_sub_fp_5_0 | l2_sub_fp_5_1;
        l3_valid_5_0 <= 1;
    end
    l3_sub_fp_5_1 <= 0;
    l3_valid_5_1  <= 0;
    if(l2_valid_5_2 | l2_valid_5_3)begin
        l3_sub_fp_5_1 <= l2_sub_fp_5_2 | l2_sub_fp_5_3;
        l3_valid_5_1 <= 1;
    end
    l3_sub_fp_5_2 <= 0;
    l3_valid_5_2  <= 0;
    if(l2_valid_5_4 | l2_valid_5_5)begin
        l3_sub_fp_5_2 <= l2_sub_fp_5_4 | l2_sub_fp_5_5;
        l3_valid_5_2 <= 1;
    end
    l3_sub_fp_5_3 <= 0;
    l3_valid_5_3  <= 0;
    if(l2_valid_5_6 | l2_valid_5_7)begin
        l3_sub_fp_5_3 <= l2_sub_fp_5_6 | l2_sub_fp_5_7;
        l3_valid_5_3 <= 1;
    end
    l3_sub_fp_6_0 <= 0;
    l3_valid_6_0  <= 0;
    if(l2_valid_6_0 | l2_valid_6_1)begin
        l3_sub_fp_6_0 <= l2_sub_fp_6_0 | l2_sub_fp_6_1;
        l3_valid_6_0 <= 1;
    end
    l3_sub_fp_6_1 <= 0;
    l3_valid_6_1  <= 0;
    if(l2_valid_6_2 | l2_valid_6_3)begin
        l3_sub_fp_6_1 <= l2_sub_fp_6_2 | l2_sub_fp_6_3;
        l3_valid_6_1 <= 1;
    end
    l3_sub_fp_6_2 <= 0;
    l3_valid_6_2  <= 0;
    if(l2_valid_6_4 | l2_valid_6_5)begin
        l3_sub_fp_6_2 <= l2_sub_fp_6_4 | l2_sub_fp_6_5;
        l3_valid_6_2 <= 1;
    end
    l3_sub_fp_6_3 <= 0;
    l3_valid_6_3  <= 0;
    if(l2_valid_6_6 | l2_valid_6_7)begin
        l3_sub_fp_6_3 <= l2_sub_fp_6_6 | l2_sub_fp_6_7;
        l3_valid_6_3 <= 1;
    end
    l3_sub_fp_7_0 <= 0;
    l3_valid_7_0  <= 0;
    if(l2_valid_7_0 | l2_valid_7_1)begin
        l3_sub_fp_7_0 <= l2_sub_fp_7_0 | l2_sub_fp_7_1;
        l3_valid_7_0 <= 1;
    end
    l3_sub_fp_7_1 <= 0;
    l3_valid_7_1  <= 0;
    if(l2_valid_7_2 | l2_valid_7_3)begin
        l3_sub_fp_7_1 <= l2_sub_fp_7_2 | l2_sub_fp_7_3;
        l3_valid_7_1 <= 1;
    end
    l3_sub_fp_7_2 <= 0;
    l3_valid_7_2  <= 0;
    if(l2_valid_7_4 | l2_valid_7_5)begin
        l3_sub_fp_7_2 <= l2_sub_fp_7_4 | l2_sub_fp_7_5;
        l3_valid_7_2 <= 1;
    end
    l3_sub_fp_7_3 <= 0;
    l3_valid_7_3  <= 0;
    if(l2_valid_7_6 | l2_valid_7_7)begin
        l3_sub_fp_7_3 <= l2_sub_fp_7_6 | l2_sub_fp_7_7;
        l3_valid_7_3 <= 1;
    end
end

//Layer 4
always@(posedge clk)begin
    l4_sub_fp_0 <= 0;
    l4_valid_0  <= 0;
    if(l3_valid_0_0 | l3_valid_0_1 |
       l3_valid_0_2 | l3_valid_0_3 )begin
        l4_sub_fp_0 <= l3_sub_fp_0_0 | l3_sub_fp_0_1 |
                          l3_sub_fp_0_2 | l3_sub_fp_0_3;
        l4_valid_0 <= 1;
    end
    l4_sub_fp_1 <= 0;
    l4_valid_1  <= 0;
    if(l3_valid_1_0 | l3_valid_1_1 |
       l3_valid_1_2 | l3_valid_1_3 )begin
        l4_sub_fp_1 <= l3_sub_fp_1_0 | l3_sub_fp_1_1 |
                          l3_sub_fp_1_2 | l3_sub_fp_1_3;
        l4_valid_1 <= 1;
    end
    l4_sub_fp_2 <= 0;
    l4_valid_2  <= 0;
    if(l3_valid_2_0 | l3_valid_2_1 |
       l3_valid_2_2 | l3_valid_2_3 )begin
        l4_sub_fp_2 <= l3_sub_fp_2_0 | l3_sub_fp_2_1 |
                          l3_sub_fp_2_2 | l3_sub_fp_2_3;
        l4_valid_2 <= 1;
    end
    l4_sub_fp_3 <= 0;
    l4_valid_3  <= 0;
    if(l3_valid_3_0 | l3_valid_3_1 |
       l3_valid_3_2 | l3_valid_3_3 )begin
        l4_sub_fp_3 <= l3_sub_fp_3_0 | l3_sub_fp_3_1 |
                          l3_sub_fp_3_2 | l3_sub_fp_3_3;
        l4_valid_3 <= 1;
    end
    l4_sub_fp_4 <= 0;
    l4_valid_4  <= 0;
    if(l3_valid_4_0 | l3_valid_4_1 |
       l3_valid_4_2 | l3_valid_4_3 )begin
        l4_sub_fp_4 <= l3_sub_fp_4_0 | l3_sub_fp_4_1 |
                          l3_sub_fp_4_2 | l3_sub_fp_4_3;
        l4_valid_4 <= 1;
    end
    l4_sub_fp_5 <= 0;
    l4_valid_5  <= 0;
    if(l3_valid_5_0 | l3_valid_5_1 |
       l3_valid_5_2 | l3_valid_5_3 )begin
        l4_sub_fp_5 <= l3_sub_fp_5_0 | l3_sub_fp_5_1 |
                          l3_sub_fp_5_2 | l3_sub_fp_5_3;
        l4_valid_5 <= 1;
    end
    l4_sub_fp_6 <= 0;
    l4_valid_6  <= 0;
    if(l3_valid_6_0 | l3_valid_6_1 |
       l3_valid_6_2 | l3_valid_6_3 )begin
        l4_sub_fp_6 <= l3_sub_fp_6_0 | l3_sub_fp_6_1 |
                          l3_sub_fp_6_2 | l3_sub_fp_6_3;
        l4_valid_6 <= 1;
    end
    l4_sub_fp_7 <= 0;
    l4_valid_7  <= 0;
    if(l3_valid_7_0 | l3_valid_7_1 |
       l3_valid_7_2 | l3_valid_7_3 )begin
        l4_sub_fp_7 <= l3_sub_fp_7_0 | l3_sub_fp_7_1 |
                          l3_sub_fp_7_2 | l3_sub_fp_7_3;
        l4_valid_7 <= 1;
    end
end

//Layer 5, accumulate
always@(posedge clk)begin
    if(rst)begin
        sub_fp_0 <= 0;
        sub_fp_1 <= 0;
        sub_fp_2 <= 0;
        sub_fp_3 <= 0;
        sub_fp_4 <= 0;
        sub_fp_5 <= 0;
        sub_fp_6 <= 0;
        sub_fp_7 <= 0;
    end else begin
        if(last_r4)begin
            sub_fp_0 <= 0;
        end else if (l4_valid_0)begin
            sub_fp_0 <= sub_fp_0 | l4_sub_fp_0;
        end
        if(last_r4)begin
            sub_fp_1 <= 0;
        end else if (l4_valid_1)begin
            sub_fp_1 <= sub_fp_1 | l4_sub_fp_1;
        end
        if(last_r4)begin
            sub_fp_2 <= 0;
        end else if (l4_valid_2)begin
            sub_fp_2 <= sub_fp_2 | l4_sub_fp_2;
        end
        if(last_r4)begin
            sub_fp_3 <= 0;
        end else if (l4_valid_3)begin
            sub_fp_3 <= sub_fp_3 | l4_sub_fp_3;
        end
        if(last_r4)begin
            sub_fp_4 <= 0;
        end else if (l4_valid_4)begin
            sub_fp_4 <= sub_fp_4 | l4_sub_fp_4;
        end
        if(last_r4)begin
            sub_fp_5 <= 0;
        end else if (l4_valid_5)begin
            sub_fp_5 <= sub_fp_5 | l4_sub_fp_5;
        end
        if(last_r4)begin
            sub_fp_6 <= 0;
        end else if (l4_valid_6)begin
            sub_fp_6 <= sub_fp_6 | l4_sub_fp_6;
        end
        if(last_r4)begin
            sub_fp_7 <= 0;
        end else if (l4_valid_7)begin
            sub_fp_7 <= sub_fp_7 | l4_sub_fp_7;
        end
    end
end


//generate fp
always@(posedge clk)begin
    if(rst)begin
        fp_valid <= 0;
        last_r1  <= 0;
        last_r2  <= 0;
        last_r3  <= 0;
        last_r4  <= 0;
    end else begin
        last_r1 <= last;
        last_r2 <= last_r1;
        last_r3 <= last_r2;
        last_r4 <= last_r3;

        fp_valid <= last_r4;
    end
    fp_data[(0+1)*BUCKET_WIDTH-1:0*BUCKET_WIDTH] <= sub_fp_0;
    fp_data[(1+1)*BUCKET_WIDTH-1:1*BUCKET_WIDTH] <= sub_fp_1;
    fp_data[(2+1)*BUCKET_WIDTH-1:2*BUCKET_WIDTH] <= sub_fp_2;
    fp_data[(3+1)*BUCKET_WIDTH-1:3*BUCKET_WIDTH] <= sub_fp_3;
    fp_data[(4+1)*BUCKET_WIDTH-1:4*BUCKET_WIDTH] <= sub_fp_4;
    fp_data[(5+1)*BUCKET_WIDTH-1:5*BUCKET_WIDTH] <= sub_fp_5;
    fp_data[(6+1)*BUCKET_WIDTH-1:6*BUCKET_WIDTH] <= sub_fp_6;
    fp_data[(7+1)*BUCKET_WIDTH-1:7*BUCKET_WIDTH] <= sub_fp_7;
end


endmodule

`include "./struct_s.sv"
module hashtable_top(clk,
	dout_0_0,dout_valid_0_0,
	dout_0_1,dout_valid_0_1,
	dout_0_2,dout_valid_0_2,
	dout_0_3,dout_valid_0_3,
	dout_0_4,dout_valid_0_4,
	dout_0_5,dout_valid_0_5,
	dout_0_6,dout_valid_0_6,
	dout_0_7,dout_valid_0_7,
	dout_0_8,dout_valid_0_8,
	dout_0_9,dout_valid_0_9,
	dout_0_10,dout_valid_0_10,
	dout_0_11,dout_valid_0_11,
	dout_0_12,dout_valid_0_12,
	dout_0_13,dout_valid_0_13,
	dout_0_14,dout_valid_0_14,
	dout_0_15,dout_valid_0_15,
	dout_0_16,dout_valid_0_16,
	dout_0_17,dout_valid_0_17,
	dout_0_18,dout_valid_0_18,
	dout_0_19,dout_valid_0_19,
	dout_0_20,dout_valid_0_20,
	dout_0_21,dout_valid_0_21,
	dout_0_22,dout_valid_0_22,
	dout_0_23,dout_valid_0_23,
	dout_0_24,dout_valid_0_24,
	dout_0_25,dout_valid_0_25,
	dout_0_26,dout_valid_0_26,
	dout_0_27,dout_valid_0_27,
	dout_0_28,dout_valid_0_28,
	dout_0_29,dout_valid_0_29,
	dout_0_30,dout_valid_0_30,
	dout_0_31,dout_valid_0_31,
	dout_1_0,dout_valid_1_0,
	dout_1_1,dout_valid_1_1,
	dout_1_2,dout_valid_1_2,
	dout_1_3,dout_valid_1_3,
	dout_1_4,dout_valid_1_4,
	dout_1_5,dout_valid_1_5,
	dout_1_6,dout_valid_1_6,
	dout_1_7,dout_valid_1_7,
	dout_1_8,dout_valid_1_8,
	dout_1_9,dout_valid_1_9,
	dout_1_10,dout_valid_1_10,
	dout_1_11,dout_valid_1_11,
	dout_1_12,dout_valid_1_12,
	dout_1_13,dout_valid_1_13,
	dout_1_14,dout_valid_1_14,
	dout_1_15,dout_valid_1_15,
	dout_1_16,dout_valid_1_16,
	dout_1_17,dout_valid_1_17,
	dout_1_18,dout_valid_1_18,
	dout_1_19,dout_valid_1_19,
	dout_1_20,dout_valid_1_20,
	dout_1_21,dout_valid_1_21,
	dout_1_22,dout_valid_1_22,
	dout_1_23,dout_valid_1_23,
	dout_1_24,dout_valid_1_24,
	dout_1_25,dout_valid_1_25,
	dout_1_26,dout_valid_1_26,
	dout_1_27,dout_valid_1_27,
	dout_1_28,dout_valid_1_28,
	dout_1_29,dout_valid_1_29,
	dout_1_30,dout_valid_1_30,
	dout_1_31,dout_valid_1_31,
	dout_2_0,dout_valid_2_0,
	dout_2_1,dout_valid_2_1,
	dout_2_2,dout_valid_2_2,
	dout_2_3,dout_valid_2_3,
	dout_2_4,dout_valid_2_4,
	dout_2_5,dout_valid_2_5,
	dout_2_6,dout_valid_2_6,
	dout_2_7,dout_valid_2_7,
	dout_2_8,dout_valid_2_8,
	dout_2_9,dout_valid_2_9,
	dout_2_10,dout_valid_2_10,
	dout_2_11,dout_valid_2_11,
	dout_2_12,dout_valid_2_12,
	dout_2_13,dout_valid_2_13,
	dout_2_14,dout_valid_2_14,
	dout_2_15,dout_valid_2_15,
	dout_2_16,dout_valid_2_16,
	dout_2_17,dout_valid_2_17,
	dout_2_18,dout_valid_2_18,
	dout_2_19,dout_valid_2_19,
	dout_2_20,dout_valid_2_20,
	dout_2_21,dout_valid_2_21,
	dout_2_22,dout_valid_2_22,
	dout_2_23,dout_valid_2_23,
	dout_2_24,dout_valid_2_24,
	dout_2_25,dout_valid_2_25,
	dout_2_26,dout_valid_2_26,
	dout_2_27,dout_valid_2_27,
	dout_2_28,dout_valid_2_28,
	dout_2_29,dout_valid_2_29,
	dout_2_30,dout_valid_2_30,
	dout_2_31,dout_valid_2_31,
	dout_3_0,dout_valid_3_0,
	dout_3_1,dout_valid_3_1,
	dout_3_2,dout_valid_3_2,
	dout_3_3,dout_valid_3_3,
	dout_3_4,dout_valid_3_4,
	dout_3_5,dout_valid_3_5,
	dout_3_6,dout_valid_3_6,
	dout_3_7,dout_valid_3_7,
	dout_3_8,dout_valid_3_8,
	dout_3_9,dout_valid_3_9,
	dout_3_10,dout_valid_3_10,
	dout_3_11,dout_valid_3_11,
	dout_3_12,dout_valid_3_12,
	dout_3_13,dout_valid_3_13,
	dout_3_14,dout_valid_3_14,
	dout_3_15,dout_valid_3_15,
	dout_3_16,dout_valid_3_16,
	dout_3_17,dout_valid_3_17,
	dout_3_18,dout_valid_3_18,
	dout_3_19,dout_valid_3_19,
	dout_3_20,dout_valid_3_20,
	dout_3_21,dout_valid_3_21,
	dout_3_22,dout_valid_3_22,
	dout_3_23,dout_valid_3_23,
	dout_3_24,dout_valid_3_24,
	dout_3_25,dout_valid_3_25,
	dout_3_26,dout_valid_3_26,
	dout_3_27,dout_valid_3_27,
	dout_3_28,dout_valid_3_28,
	dout_3_29,dout_valid_3_29,
	dout_3_30,dout_valid_3_30,
	dout_3_31,dout_valid_3_31,
	dout_4_0,dout_valid_4_0,
	dout_4_1,dout_valid_4_1,
	dout_4_2,dout_valid_4_2,
	dout_4_3,dout_valid_4_3,
	dout_4_4,dout_valid_4_4,
	dout_4_5,dout_valid_4_5,
	dout_4_6,dout_valid_4_6,
	dout_4_7,dout_valid_4_7,
	dout_4_8,dout_valid_4_8,
	dout_4_9,dout_valid_4_9,
	dout_4_10,dout_valid_4_10,
	dout_4_11,dout_valid_4_11,
	dout_4_12,dout_valid_4_12,
	dout_4_13,dout_valid_4_13,
	dout_4_14,dout_valid_4_14,
	dout_4_15,dout_valid_4_15,
	dout_4_16,dout_valid_4_16,
	dout_4_17,dout_valid_4_17,
	dout_4_18,dout_valid_4_18,
	dout_4_19,dout_valid_4_19,
	dout_4_20,dout_valid_4_20,
	dout_4_21,dout_valid_4_21,
	dout_4_22,dout_valid_4_22,
	dout_4_23,dout_valid_4_23,
	dout_4_24,dout_valid_4_24,
	dout_4_25,dout_valid_4_25,
	dout_4_26,dout_valid_4_26,
	dout_4_27,dout_valid_4_27,
	dout_4_28,dout_valid_4_28,
	dout_4_29,dout_valid_4_29,
	dout_4_30,dout_valid_4_30,
	dout_4_31,dout_valid_4_31,
	dout_5_0,dout_valid_5_0,
	dout_5_1,dout_valid_5_1,
	dout_5_2,dout_valid_5_2,
	dout_5_3,dout_valid_5_3,
	dout_5_4,dout_valid_5_4,
	dout_5_5,dout_valid_5_5,
	dout_5_6,dout_valid_5_6,
	dout_5_7,dout_valid_5_7,
	dout_5_8,dout_valid_5_8,
	dout_5_9,dout_valid_5_9,
	dout_5_10,dout_valid_5_10,
	dout_5_11,dout_valid_5_11,
	dout_5_12,dout_valid_5_12,
	dout_5_13,dout_valid_5_13,
	dout_5_14,dout_valid_5_14,
	dout_5_15,dout_valid_5_15,
	dout_5_16,dout_valid_5_16,
	dout_5_17,dout_valid_5_17,
	dout_5_18,dout_valid_5_18,
	dout_5_19,dout_valid_5_19,
	dout_5_20,dout_valid_5_20,
	dout_5_21,dout_valid_5_21,
	dout_5_22,dout_valid_5_22,
	dout_5_23,dout_valid_5_23,
	dout_5_24,dout_valid_5_24,
	dout_5_25,dout_valid_5_25,
	dout_5_26,dout_valid_5_26,
	dout_5_27,dout_valid_5_27,
	dout_5_28,dout_valid_5_28,
	dout_5_29,dout_valid_5_29,
	dout_5_30,dout_valid_5_30,
	dout_5_31,dout_valid_5_31,
	dout_6_0,dout_valid_6_0,
	dout_6_1,dout_valid_6_1,
	dout_6_2,dout_valid_6_2,
	dout_6_3,dout_valid_6_3,
	dout_6_4,dout_valid_6_4,
	dout_6_5,dout_valid_6_5,
	dout_6_6,dout_valid_6_6,
	dout_6_7,dout_valid_6_7,
	dout_6_8,dout_valid_6_8,
	dout_6_9,dout_valid_6_9,
	dout_6_10,dout_valid_6_10,
	dout_6_11,dout_valid_6_11,
	dout_6_12,dout_valid_6_12,
	dout_6_13,dout_valid_6_13,
	dout_6_14,dout_valid_6_14,
	dout_6_15,dout_valid_6_15,
	dout_6_16,dout_valid_6_16,
	dout_6_17,dout_valid_6_17,
	dout_6_18,dout_valid_6_18,
	dout_6_19,dout_valid_6_19,
	dout_6_20,dout_valid_6_20,
	dout_6_21,dout_valid_6_21,
	dout_6_22,dout_valid_6_22,
	dout_6_23,dout_valid_6_23,
	dout_6_24,dout_valid_6_24,
	dout_6_25,dout_valid_6_25,
	dout_6_26,dout_valid_6_26,
	dout_6_27,dout_valid_6_27,
	dout_6_28,dout_valid_6_28,
	dout_6_29,dout_valid_6_29,
	dout_6_30,dout_valid_6_30,
	dout_6_31,dout_valid_6_31,
	dout_7_0,dout_valid_7_0,
	dout_7_1,dout_valid_7_1,
	dout_7_2,dout_valid_7_2,
	dout_7_3,dout_valid_7_3,
	dout_7_4,dout_valid_7_4,
	dout_7_5,dout_valid_7_5,
	dout_7_6,dout_valid_7_6,
	dout_7_7,dout_valid_7_7,
	dout_7_8,dout_valid_7_8,
	dout_7_9,dout_valid_7_9,
	dout_7_10,dout_valid_7_10,
	dout_7_11,dout_valid_7_11,
	dout_7_12,dout_valid_7_12,
	dout_7_13,dout_valid_7_13,
	dout_7_14,dout_valid_7_14,
	dout_7_15,dout_valid_7_15,
	dout_7_16,dout_valid_7_16,
	dout_7_17,dout_valid_7_17,
	dout_7_18,dout_valid_7_18,
	dout_7_19,dout_valid_7_19,
	dout_7_20,dout_valid_7_20,
	dout_7_21,dout_valid_7_21,
	dout_7_22,dout_valid_7_22,
	dout_7_23,dout_valid_7_23,
	dout_7_24,dout_valid_7_24,
	dout_7_25,dout_valid_7_25,
	dout_7_26,dout_valid_7_26,
	dout_7_27,dout_valid_7_27,
	dout_7_28,dout_valid_7_28,
	dout_7_29,dout_valid_7_29,
	dout_7_30,dout_valid_7_30,
	dout_7_31,dout_valid_7_31,
    din,din_valid
);

input clk;
input [255:0] din;
input din_valid;
output wire [RID_WIDTH-1:0] dout_0_0;
output wire dout_valid_0_0;
output wire [RID_WIDTH-1:0] dout_0_1;
output wire dout_valid_0_1;
output wire [RID_WIDTH-1:0] dout_0_2;
output wire dout_valid_0_2;
output wire [RID_WIDTH-1:0] dout_0_3;
output wire dout_valid_0_3;
output wire [RID_WIDTH-1:0] dout_0_4;
output wire dout_valid_0_4;
output wire [RID_WIDTH-1:0] dout_0_5;
output wire dout_valid_0_5;
output wire [RID_WIDTH-1:0] dout_0_6;
output wire dout_valid_0_6;
output wire [RID_WIDTH-1:0] dout_0_7;
output wire dout_valid_0_7;
output wire [RID_WIDTH-1:0] dout_0_8;
output wire dout_valid_0_8;
output wire [RID_WIDTH-1:0] dout_0_9;
output wire dout_valid_0_9;
output wire [RID_WIDTH-1:0] dout_0_10;
output wire dout_valid_0_10;
output wire [RID_WIDTH-1:0] dout_0_11;
output wire dout_valid_0_11;
output wire [RID_WIDTH-1:0] dout_0_12;
output wire dout_valid_0_12;
output wire [RID_WIDTH-1:0] dout_0_13;
output wire dout_valid_0_13;
output wire [RID_WIDTH-1:0] dout_0_14;
output wire dout_valid_0_14;
output wire [RID_WIDTH-1:0] dout_0_15;
output wire dout_valid_0_15;
output wire [RID_WIDTH-1:0] dout_0_16;
output wire dout_valid_0_16;
output wire [RID_WIDTH-1:0] dout_0_17;
output wire dout_valid_0_17;
output wire [RID_WIDTH-1:0] dout_0_18;
output wire dout_valid_0_18;
output wire [RID_WIDTH-1:0] dout_0_19;
output wire dout_valid_0_19;
output wire [RID_WIDTH-1:0] dout_0_20;
output wire dout_valid_0_20;
output wire [RID_WIDTH-1:0] dout_0_21;
output wire dout_valid_0_21;
output wire [RID_WIDTH-1:0] dout_0_22;
output wire dout_valid_0_22;
output wire [RID_WIDTH-1:0] dout_0_23;
output wire dout_valid_0_23;
output wire [RID_WIDTH-1:0] dout_0_24;
output wire dout_valid_0_24;
output wire [RID_WIDTH-1:0] dout_0_25;
output wire dout_valid_0_25;
output wire [RID_WIDTH-1:0] dout_0_26;
output wire dout_valid_0_26;
output wire [RID_WIDTH-1:0] dout_0_27;
output wire dout_valid_0_27;
output wire [RID_WIDTH-1:0] dout_0_28;
output wire dout_valid_0_28;
output wire [RID_WIDTH-1:0] dout_0_29;
output wire dout_valid_0_29;
output wire [RID_WIDTH-1:0] dout_0_30;
output wire dout_valid_0_30;
output wire [RID_WIDTH-1:0] dout_0_31;
output wire dout_valid_0_31;
output wire [RID_WIDTH-1:0] dout_1_0;
output wire dout_valid_1_0;
output wire [RID_WIDTH-1:0] dout_1_1;
output wire dout_valid_1_1;
output wire [RID_WIDTH-1:0] dout_1_2;
output wire dout_valid_1_2;
output wire [RID_WIDTH-1:0] dout_1_3;
output wire dout_valid_1_3;
output wire [RID_WIDTH-1:0] dout_1_4;
output wire dout_valid_1_4;
output wire [RID_WIDTH-1:0] dout_1_5;
output wire dout_valid_1_5;
output wire [RID_WIDTH-1:0] dout_1_6;
output wire dout_valid_1_6;
output wire [RID_WIDTH-1:0] dout_1_7;
output wire dout_valid_1_7;
output wire [RID_WIDTH-1:0] dout_1_8;
output wire dout_valid_1_8;
output wire [RID_WIDTH-1:0] dout_1_9;
output wire dout_valid_1_9;
output wire [RID_WIDTH-1:0] dout_1_10;
output wire dout_valid_1_10;
output wire [RID_WIDTH-1:0] dout_1_11;
output wire dout_valid_1_11;
output wire [RID_WIDTH-1:0] dout_1_12;
output wire dout_valid_1_12;
output wire [RID_WIDTH-1:0] dout_1_13;
output wire dout_valid_1_13;
output wire [RID_WIDTH-1:0] dout_1_14;
output wire dout_valid_1_14;
output wire [RID_WIDTH-1:0] dout_1_15;
output wire dout_valid_1_15;
output wire [RID_WIDTH-1:0] dout_1_16;
output wire dout_valid_1_16;
output wire [RID_WIDTH-1:0] dout_1_17;
output wire dout_valid_1_17;
output wire [RID_WIDTH-1:0] dout_1_18;
output wire dout_valid_1_18;
output wire [RID_WIDTH-1:0] dout_1_19;
output wire dout_valid_1_19;
output wire [RID_WIDTH-1:0] dout_1_20;
output wire dout_valid_1_20;
output wire [RID_WIDTH-1:0] dout_1_21;
output wire dout_valid_1_21;
output wire [RID_WIDTH-1:0] dout_1_22;
output wire dout_valid_1_22;
output wire [RID_WIDTH-1:0] dout_1_23;
output wire dout_valid_1_23;
output wire [RID_WIDTH-1:0] dout_1_24;
output wire dout_valid_1_24;
output wire [RID_WIDTH-1:0] dout_1_25;
output wire dout_valid_1_25;
output wire [RID_WIDTH-1:0] dout_1_26;
output wire dout_valid_1_26;
output wire [RID_WIDTH-1:0] dout_1_27;
output wire dout_valid_1_27;
output wire [RID_WIDTH-1:0] dout_1_28;
output wire dout_valid_1_28;
output wire [RID_WIDTH-1:0] dout_1_29;
output wire dout_valid_1_29;
output wire [RID_WIDTH-1:0] dout_1_30;
output wire dout_valid_1_30;
output wire [RID_WIDTH-1:0] dout_1_31;
output wire dout_valid_1_31;
output wire [RID_WIDTH-1:0] dout_2_0;
output wire dout_valid_2_0;
output wire [RID_WIDTH-1:0] dout_2_1;
output wire dout_valid_2_1;
output wire [RID_WIDTH-1:0] dout_2_2;
output wire dout_valid_2_2;
output wire [RID_WIDTH-1:0] dout_2_3;
output wire dout_valid_2_3;
output wire [RID_WIDTH-1:0] dout_2_4;
output wire dout_valid_2_4;
output wire [RID_WIDTH-1:0] dout_2_5;
output wire dout_valid_2_5;
output wire [RID_WIDTH-1:0] dout_2_6;
output wire dout_valid_2_6;
output wire [RID_WIDTH-1:0] dout_2_7;
output wire dout_valid_2_7;
output wire [RID_WIDTH-1:0] dout_2_8;
output wire dout_valid_2_8;
output wire [RID_WIDTH-1:0] dout_2_9;
output wire dout_valid_2_9;
output wire [RID_WIDTH-1:0] dout_2_10;
output wire dout_valid_2_10;
output wire [RID_WIDTH-1:0] dout_2_11;
output wire dout_valid_2_11;
output wire [RID_WIDTH-1:0] dout_2_12;
output wire dout_valid_2_12;
output wire [RID_WIDTH-1:0] dout_2_13;
output wire dout_valid_2_13;
output wire [RID_WIDTH-1:0] dout_2_14;
output wire dout_valid_2_14;
output wire [RID_WIDTH-1:0] dout_2_15;
output wire dout_valid_2_15;
output wire [RID_WIDTH-1:0] dout_2_16;
output wire dout_valid_2_16;
output wire [RID_WIDTH-1:0] dout_2_17;
output wire dout_valid_2_17;
output wire [RID_WIDTH-1:0] dout_2_18;
output wire dout_valid_2_18;
output wire [RID_WIDTH-1:0] dout_2_19;
output wire dout_valid_2_19;
output wire [RID_WIDTH-1:0] dout_2_20;
output wire dout_valid_2_20;
output wire [RID_WIDTH-1:0] dout_2_21;
output wire dout_valid_2_21;
output wire [RID_WIDTH-1:0] dout_2_22;
output wire dout_valid_2_22;
output wire [RID_WIDTH-1:0] dout_2_23;
output wire dout_valid_2_23;
output wire [RID_WIDTH-1:0] dout_2_24;
output wire dout_valid_2_24;
output wire [RID_WIDTH-1:0] dout_2_25;
output wire dout_valid_2_25;
output wire [RID_WIDTH-1:0] dout_2_26;
output wire dout_valid_2_26;
output wire [RID_WIDTH-1:0] dout_2_27;
output wire dout_valid_2_27;
output wire [RID_WIDTH-1:0] dout_2_28;
output wire dout_valid_2_28;
output wire [RID_WIDTH-1:0] dout_2_29;
output wire dout_valid_2_29;
output wire [RID_WIDTH-1:0] dout_2_30;
output wire dout_valid_2_30;
output wire [RID_WIDTH-1:0] dout_2_31;
output wire dout_valid_2_31;
output wire [RID_WIDTH-1:0] dout_3_0;
output wire dout_valid_3_0;
output wire [RID_WIDTH-1:0] dout_3_1;
output wire dout_valid_3_1;
output wire [RID_WIDTH-1:0] dout_3_2;
output wire dout_valid_3_2;
output wire [RID_WIDTH-1:0] dout_3_3;
output wire dout_valid_3_3;
output wire [RID_WIDTH-1:0] dout_3_4;
output wire dout_valid_3_4;
output wire [RID_WIDTH-1:0] dout_3_5;
output wire dout_valid_3_5;
output wire [RID_WIDTH-1:0] dout_3_6;
output wire dout_valid_3_6;
output wire [RID_WIDTH-1:0] dout_3_7;
output wire dout_valid_3_7;
output wire [RID_WIDTH-1:0] dout_3_8;
output wire dout_valid_3_8;
output wire [RID_WIDTH-1:0] dout_3_9;
output wire dout_valid_3_9;
output wire [RID_WIDTH-1:0] dout_3_10;
output wire dout_valid_3_10;
output wire [RID_WIDTH-1:0] dout_3_11;
output wire dout_valid_3_11;
output wire [RID_WIDTH-1:0] dout_3_12;
output wire dout_valid_3_12;
output wire [RID_WIDTH-1:0] dout_3_13;
output wire dout_valid_3_13;
output wire [RID_WIDTH-1:0] dout_3_14;
output wire dout_valid_3_14;
output wire [RID_WIDTH-1:0] dout_3_15;
output wire dout_valid_3_15;
output wire [RID_WIDTH-1:0] dout_3_16;
output wire dout_valid_3_16;
output wire [RID_WIDTH-1:0] dout_3_17;
output wire dout_valid_3_17;
output wire [RID_WIDTH-1:0] dout_3_18;
output wire dout_valid_3_18;
output wire [RID_WIDTH-1:0] dout_3_19;
output wire dout_valid_3_19;
output wire [RID_WIDTH-1:0] dout_3_20;
output wire dout_valid_3_20;
output wire [RID_WIDTH-1:0] dout_3_21;
output wire dout_valid_3_21;
output wire [RID_WIDTH-1:0] dout_3_22;
output wire dout_valid_3_22;
output wire [RID_WIDTH-1:0] dout_3_23;
output wire dout_valid_3_23;
output wire [RID_WIDTH-1:0] dout_3_24;
output wire dout_valid_3_24;
output wire [RID_WIDTH-1:0] dout_3_25;
output wire dout_valid_3_25;
output wire [RID_WIDTH-1:0] dout_3_26;
output wire dout_valid_3_26;
output wire [RID_WIDTH-1:0] dout_3_27;
output wire dout_valid_3_27;
output wire [RID_WIDTH-1:0] dout_3_28;
output wire dout_valid_3_28;
output wire [RID_WIDTH-1:0] dout_3_29;
output wire dout_valid_3_29;
output wire [RID_WIDTH-1:0] dout_3_30;
output wire dout_valid_3_30;
output wire [RID_WIDTH-1:0] dout_3_31;
output wire dout_valid_3_31;
output wire [RID_WIDTH-1:0] dout_4_0;
output wire dout_valid_4_0;
output wire [RID_WIDTH-1:0] dout_4_1;
output wire dout_valid_4_1;
output wire [RID_WIDTH-1:0] dout_4_2;
output wire dout_valid_4_2;
output wire [RID_WIDTH-1:0] dout_4_3;
output wire dout_valid_4_3;
output wire [RID_WIDTH-1:0] dout_4_4;
output wire dout_valid_4_4;
output wire [RID_WIDTH-1:0] dout_4_5;
output wire dout_valid_4_5;
output wire [RID_WIDTH-1:0] dout_4_6;
output wire dout_valid_4_6;
output wire [RID_WIDTH-1:0] dout_4_7;
output wire dout_valid_4_7;
output wire [RID_WIDTH-1:0] dout_4_8;
output wire dout_valid_4_8;
output wire [RID_WIDTH-1:0] dout_4_9;
output wire dout_valid_4_9;
output wire [RID_WIDTH-1:0] dout_4_10;
output wire dout_valid_4_10;
output wire [RID_WIDTH-1:0] dout_4_11;
output wire dout_valid_4_11;
output wire [RID_WIDTH-1:0] dout_4_12;
output wire dout_valid_4_12;
output wire [RID_WIDTH-1:0] dout_4_13;
output wire dout_valid_4_13;
output wire [RID_WIDTH-1:0] dout_4_14;
output wire dout_valid_4_14;
output wire [RID_WIDTH-1:0] dout_4_15;
output wire dout_valid_4_15;
output wire [RID_WIDTH-1:0] dout_4_16;
output wire dout_valid_4_16;
output wire [RID_WIDTH-1:0] dout_4_17;
output wire dout_valid_4_17;
output wire [RID_WIDTH-1:0] dout_4_18;
output wire dout_valid_4_18;
output wire [RID_WIDTH-1:0] dout_4_19;
output wire dout_valid_4_19;
output wire [RID_WIDTH-1:0] dout_4_20;
output wire dout_valid_4_20;
output wire [RID_WIDTH-1:0] dout_4_21;
output wire dout_valid_4_21;
output wire [RID_WIDTH-1:0] dout_4_22;
output wire dout_valid_4_22;
output wire [RID_WIDTH-1:0] dout_4_23;
output wire dout_valid_4_23;
output wire [RID_WIDTH-1:0] dout_4_24;
output wire dout_valid_4_24;
output wire [RID_WIDTH-1:0] dout_4_25;
output wire dout_valid_4_25;
output wire [RID_WIDTH-1:0] dout_4_26;
output wire dout_valid_4_26;
output wire [RID_WIDTH-1:0] dout_4_27;
output wire dout_valid_4_27;
output wire [RID_WIDTH-1:0] dout_4_28;
output wire dout_valid_4_28;
output wire [RID_WIDTH-1:0] dout_4_29;
output wire dout_valid_4_29;
output wire [RID_WIDTH-1:0] dout_4_30;
output wire dout_valid_4_30;
output wire [RID_WIDTH-1:0] dout_4_31;
output wire dout_valid_4_31;
output wire [RID_WIDTH-1:0] dout_5_0;
output wire dout_valid_5_0;
output wire [RID_WIDTH-1:0] dout_5_1;
output wire dout_valid_5_1;
output wire [RID_WIDTH-1:0] dout_5_2;
output wire dout_valid_5_2;
output wire [RID_WIDTH-1:0] dout_5_3;
output wire dout_valid_5_3;
output wire [RID_WIDTH-1:0] dout_5_4;
output wire dout_valid_5_4;
output wire [RID_WIDTH-1:0] dout_5_5;
output wire dout_valid_5_5;
output wire [RID_WIDTH-1:0] dout_5_6;
output wire dout_valid_5_6;
output wire [RID_WIDTH-1:0] dout_5_7;
output wire dout_valid_5_7;
output wire [RID_WIDTH-1:0] dout_5_8;
output wire dout_valid_5_8;
output wire [RID_WIDTH-1:0] dout_5_9;
output wire dout_valid_5_9;
output wire [RID_WIDTH-1:0] dout_5_10;
output wire dout_valid_5_10;
output wire [RID_WIDTH-1:0] dout_5_11;
output wire dout_valid_5_11;
output wire [RID_WIDTH-1:0] dout_5_12;
output wire dout_valid_5_12;
output wire [RID_WIDTH-1:0] dout_5_13;
output wire dout_valid_5_13;
output wire [RID_WIDTH-1:0] dout_5_14;
output wire dout_valid_5_14;
output wire [RID_WIDTH-1:0] dout_5_15;
output wire dout_valid_5_15;
output wire [RID_WIDTH-1:0] dout_5_16;
output wire dout_valid_5_16;
output wire [RID_WIDTH-1:0] dout_5_17;
output wire dout_valid_5_17;
output wire [RID_WIDTH-1:0] dout_5_18;
output wire dout_valid_5_18;
output wire [RID_WIDTH-1:0] dout_5_19;
output wire dout_valid_5_19;
output wire [RID_WIDTH-1:0] dout_5_20;
output wire dout_valid_5_20;
output wire [RID_WIDTH-1:0] dout_5_21;
output wire dout_valid_5_21;
output wire [RID_WIDTH-1:0] dout_5_22;
output wire dout_valid_5_22;
output wire [RID_WIDTH-1:0] dout_5_23;
output wire dout_valid_5_23;
output wire [RID_WIDTH-1:0] dout_5_24;
output wire dout_valid_5_24;
output wire [RID_WIDTH-1:0] dout_5_25;
output wire dout_valid_5_25;
output wire [RID_WIDTH-1:0] dout_5_26;
output wire dout_valid_5_26;
output wire [RID_WIDTH-1:0] dout_5_27;
output wire dout_valid_5_27;
output wire [RID_WIDTH-1:0] dout_5_28;
output wire dout_valid_5_28;
output wire [RID_WIDTH-1:0] dout_5_29;
output wire dout_valid_5_29;
output wire [RID_WIDTH-1:0] dout_5_30;
output wire dout_valid_5_30;
output wire [RID_WIDTH-1:0] dout_5_31;
output wire dout_valid_5_31;
output wire [RID_WIDTH-1:0] dout_6_0;
output wire dout_valid_6_0;
output wire [RID_WIDTH-1:0] dout_6_1;
output wire dout_valid_6_1;
output wire [RID_WIDTH-1:0] dout_6_2;
output wire dout_valid_6_2;
output wire [RID_WIDTH-1:0] dout_6_3;
output wire dout_valid_6_3;
output wire [RID_WIDTH-1:0] dout_6_4;
output wire dout_valid_6_4;
output wire [RID_WIDTH-1:0] dout_6_5;
output wire dout_valid_6_5;
output wire [RID_WIDTH-1:0] dout_6_6;
output wire dout_valid_6_6;
output wire [RID_WIDTH-1:0] dout_6_7;
output wire dout_valid_6_7;
output wire [RID_WIDTH-1:0] dout_6_8;
output wire dout_valid_6_8;
output wire [RID_WIDTH-1:0] dout_6_9;
output wire dout_valid_6_9;
output wire [RID_WIDTH-1:0] dout_6_10;
output wire dout_valid_6_10;
output wire [RID_WIDTH-1:0] dout_6_11;
output wire dout_valid_6_11;
output wire [RID_WIDTH-1:0] dout_6_12;
output wire dout_valid_6_12;
output wire [RID_WIDTH-1:0] dout_6_13;
output wire dout_valid_6_13;
output wire [RID_WIDTH-1:0] dout_6_14;
output wire dout_valid_6_14;
output wire [RID_WIDTH-1:0] dout_6_15;
output wire dout_valid_6_15;
output wire [RID_WIDTH-1:0] dout_6_16;
output wire dout_valid_6_16;
output wire [RID_WIDTH-1:0] dout_6_17;
output wire dout_valid_6_17;
output wire [RID_WIDTH-1:0] dout_6_18;
output wire dout_valid_6_18;
output wire [RID_WIDTH-1:0] dout_6_19;
output wire dout_valid_6_19;
output wire [RID_WIDTH-1:0] dout_6_20;
output wire dout_valid_6_20;
output wire [RID_WIDTH-1:0] dout_6_21;
output wire dout_valid_6_21;
output wire [RID_WIDTH-1:0] dout_6_22;
output wire dout_valid_6_22;
output wire [RID_WIDTH-1:0] dout_6_23;
output wire dout_valid_6_23;
output wire [RID_WIDTH-1:0] dout_6_24;
output wire dout_valid_6_24;
output wire [RID_WIDTH-1:0] dout_6_25;
output wire dout_valid_6_25;
output wire [RID_WIDTH-1:0] dout_6_26;
output wire dout_valid_6_26;
output wire [RID_WIDTH-1:0] dout_6_27;
output wire dout_valid_6_27;
output wire [RID_WIDTH-1:0] dout_6_28;
output wire dout_valid_6_28;
output wire [RID_WIDTH-1:0] dout_6_29;
output wire dout_valid_6_29;
output wire [RID_WIDTH-1:0] dout_6_30;
output wire dout_valid_6_30;
output wire [RID_WIDTH-1:0] dout_6_31;
output wire dout_valid_6_31;
output wire [RID_WIDTH-1:0] dout_7_0;
output wire dout_valid_7_0;
output wire [RID_WIDTH-1:0] dout_7_1;
output wire dout_valid_7_1;
output wire [RID_WIDTH-1:0] dout_7_2;
output wire dout_valid_7_2;
output wire [RID_WIDTH-1:0] dout_7_3;
output wire dout_valid_7_3;
output wire [RID_WIDTH-1:0] dout_7_4;
output wire dout_valid_7_4;
output wire [RID_WIDTH-1:0] dout_7_5;
output wire dout_valid_7_5;
output wire [RID_WIDTH-1:0] dout_7_6;
output wire dout_valid_7_6;
output wire [RID_WIDTH-1:0] dout_7_7;
output wire dout_valid_7_7;
output wire [RID_WIDTH-1:0] dout_7_8;
output wire dout_valid_7_8;
output wire [RID_WIDTH-1:0] dout_7_9;
output wire dout_valid_7_9;
output wire [RID_WIDTH-1:0] dout_7_10;
output wire dout_valid_7_10;
output wire [RID_WIDTH-1:0] dout_7_11;
output wire dout_valid_7_11;
output wire [RID_WIDTH-1:0] dout_7_12;
output wire dout_valid_7_12;
output wire [RID_WIDTH-1:0] dout_7_13;
output wire dout_valid_7_13;
output wire [RID_WIDTH-1:0] dout_7_14;
output wire dout_valid_7_14;
output wire [RID_WIDTH-1:0] dout_7_15;
output wire dout_valid_7_15;
output wire [RID_WIDTH-1:0] dout_7_16;
output wire dout_valid_7_16;
output wire [RID_WIDTH-1:0] dout_7_17;
output wire dout_valid_7_17;
output wire [RID_WIDTH-1:0] dout_7_18;
output wire dout_valid_7_18;
output wire [RID_WIDTH-1:0] dout_7_19;
output wire dout_valid_7_19;
output wire [RID_WIDTH-1:0] dout_7_20;
output wire dout_valid_7_20;
output wire [RID_WIDTH-1:0] dout_7_21;
output wire dout_valid_7_21;
output wire [RID_WIDTH-1:0] dout_7_22;
output wire dout_valid_7_22;
output wire [RID_WIDTH-1:0] dout_7_23;
output wire dout_valid_7_23;
output wire [RID_WIDTH-1:0] dout_7_24;
output wire dout_valid_7_24;
output wire [RID_WIDTH-1:0] dout_7_25;
output wire dout_valid_7_25;
output wire [RID_WIDTH-1:0] dout_7_26;
output wire dout_valid_7_26;
output wire [RID_WIDTH-1:0] dout_7_27;
output wire dout_valid_7_27;
output wire [RID_WIDTH-1:0] dout_7_28;
output wire dout_valid_7_28;
output wire [RID_WIDTH-1:0] dout_7_29;
output wire dout_valid_7_29;
output wire [RID_WIDTH-1:0] dout_7_30;
output wire dout_valid_7_30;
output wire [RID_WIDTH-1:0] dout_7_31;
output wire dout_valid_7_31;

wire [63:0] din_0_0;
wire din_valid_0_0;
wire [63:0] din_0_1;
wire din_valid_0_1;
wire [63:0] din_0_2;
wire din_valid_0_2;
wire [63:0] din_0_3;
wire din_valid_0_3;
wire [63:0] din_0_4;
wire din_valid_0_4;
wire [63:0] din_0_5;
wire din_valid_0_5;
wire [63:0] din_0_6;
wire din_valid_0_6;
wire [63:0] din_0_7;
wire din_valid_0_7;
wire [63:0] din_0_8;
wire din_valid_0_8;
wire [63:0] din_0_9;
wire din_valid_0_9;
wire [63:0] din_0_10;
wire din_valid_0_10;
wire [63:0] din_0_11;
wire din_valid_0_11;
wire [63:0] din_0_12;
wire din_valid_0_12;
wire [63:0] din_0_13;
wire din_valid_0_13;
wire [63:0] din_0_14;
wire din_valid_0_14;
wire [63:0] din_0_15;
wire din_valid_0_15;
wire [63:0] din_0_16;
wire din_valid_0_16;
wire [63:0] din_0_17;
wire din_valid_0_17;
wire [63:0] din_0_18;
wire din_valid_0_18;
wire [63:0] din_0_19;
wire din_valid_0_19;
wire [63:0] din_0_20;
wire din_valid_0_20;
wire [63:0] din_0_21;
wire din_valid_0_21;
wire [63:0] din_0_22;
wire din_valid_0_22;
wire [63:0] din_0_23;
wire din_valid_0_23;
wire [63:0] din_0_24;
wire din_valid_0_24;
wire [63:0] din_0_25;
wire din_valid_0_25;
wire [63:0] din_0_26;
wire din_valid_0_26;
wire [63:0] din_0_27;
wire din_valid_0_27;
wire [63:0] din_0_28;
wire din_valid_0_28;
wire [63:0] din_0_29;
wire din_valid_0_29;
wire [63:0] din_0_30;
wire din_valid_0_30;
wire [63:0] din_0_31;
wire din_valid_0_31;
wire [63:0] din_1_0;
wire din_valid_1_0;
wire [63:0] din_1_1;
wire din_valid_1_1;
wire [63:0] din_1_2;
wire din_valid_1_2;
wire [63:0] din_1_3;
wire din_valid_1_3;
wire [63:0] din_1_4;
wire din_valid_1_4;
wire [63:0] din_1_5;
wire din_valid_1_5;
wire [63:0] din_1_6;
wire din_valid_1_6;
wire [63:0] din_1_7;
wire din_valid_1_7;
wire [63:0] din_1_8;
wire din_valid_1_8;
wire [63:0] din_1_9;
wire din_valid_1_9;
wire [63:0] din_1_10;
wire din_valid_1_10;
wire [63:0] din_1_11;
wire din_valid_1_11;
wire [63:0] din_1_12;
wire din_valid_1_12;
wire [63:0] din_1_13;
wire din_valid_1_13;
wire [63:0] din_1_14;
wire din_valid_1_14;
wire [63:0] din_1_15;
wire din_valid_1_15;
wire [63:0] din_1_16;
wire din_valid_1_16;
wire [63:0] din_1_17;
wire din_valid_1_17;
wire [63:0] din_1_18;
wire din_valid_1_18;
wire [63:0] din_1_19;
wire din_valid_1_19;
wire [63:0] din_1_20;
wire din_valid_1_20;
wire [63:0] din_1_21;
wire din_valid_1_21;
wire [63:0] din_1_22;
wire din_valid_1_22;
wire [63:0] din_1_23;
wire din_valid_1_23;
wire [63:0] din_1_24;
wire din_valid_1_24;
wire [63:0] din_1_25;
wire din_valid_1_25;
wire [63:0] din_1_26;
wire din_valid_1_26;
wire [63:0] din_1_27;
wire din_valid_1_27;
wire [63:0] din_1_28;
wire din_valid_1_28;
wire [63:0] din_1_29;
wire din_valid_1_29;
wire [63:0] din_1_30;
wire din_valid_1_30;
wire [63:0] din_1_31;
wire din_valid_1_31;
wire [63:0] din_2_0;
wire din_valid_2_0;
wire [63:0] din_2_1;
wire din_valid_2_1;
wire [63:0] din_2_2;
wire din_valid_2_2;
wire [63:0] din_2_3;
wire din_valid_2_3;
wire [63:0] din_2_4;
wire din_valid_2_4;
wire [63:0] din_2_5;
wire din_valid_2_5;
wire [63:0] din_2_6;
wire din_valid_2_6;
wire [63:0] din_2_7;
wire din_valid_2_7;
wire [63:0] din_2_8;
wire din_valid_2_8;
wire [63:0] din_2_9;
wire din_valid_2_9;
wire [63:0] din_2_10;
wire din_valid_2_10;
wire [63:0] din_2_11;
wire din_valid_2_11;
wire [63:0] din_2_12;
wire din_valid_2_12;
wire [63:0] din_2_13;
wire din_valid_2_13;
wire [63:0] din_2_14;
wire din_valid_2_14;
wire [63:0] din_2_15;
wire din_valid_2_15;
wire [63:0] din_2_16;
wire din_valid_2_16;
wire [63:0] din_2_17;
wire din_valid_2_17;
wire [63:0] din_2_18;
wire din_valid_2_18;
wire [63:0] din_2_19;
wire din_valid_2_19;
wire [63:0] din_2_20;
wire din_valid_2_20;
wire [63:0] din_2_21;
wire din_valid_2_21;
wire [63:0] din_2_22;
wire din_valid_2_22;
wire [63:0] din_2_23;
wire din_valid_2_23;
wire [63:0] din_2_24;
wire din_valid_2_24;
wire [63:0] din_2_25;
wire din_valid_2_25;
wire [63:0] din_2_26;
wire din_valid_2_26;
wire [63:0] din_2_27;
wire din_valid_2_27;
wire [63:0] din_2_28;
wire din_valid_2_28;
wire [63:0] din_2_29;
wire din_valid_2_29;
wire [63:0] din_2_30;
wire din_valid_2_30;
wire [63:0] din_2_31;
wire din_valid_2_31;
wire [63:0] din_3_0;
wire din_valid_3_0;
wire [63:0] din_3_1;
wire din_valid_3_1;
wire [63:0] din_3_2;
wire din_valid_3_2;
wire [63:0] din_3_3;
wire din_valid_3_3;
wire [63:0] din_3_4;
wire din_valid_3_4;
wire [63:0] din_3_5;
wire din_valid_3_5;
wire [63:0] din_3_6;
wire din_valid_3_6;
wire [63:0] din_3_7;
wire din_valid_3_7;
wire [63:0] din_3_8;
wire din_valid_3_8;
wire [63:0] din_3_9;
wire din_valid_3_9;
wire [63:0] din_3_10;
wire din_valid_3_10;
wire [63:0] din_3_11;
wire din_valid_3_11;
wire [63:0] din_3_12;
wire din_valid_3_12;
wire [63:0] din_3_13;
wire din_valid_3_13;
wire [63:0] din_3_14;
wire din_valid_3_14;
wire [63:0] din_3_15;
wire din_valid_3_15;
wire [63:0] din_3_16;
wire din_valid_3_16;
wire [63:0] din_3_17;
wire din_valid_3_17;
wire [63:0] din_3_18;
wire din_valid_3_18;
wire [63:0] din_3_19;
wire din_valid_3_19;
wire [63:0] din_3_20;
wire din_valid_3_20;
wire [63:0] din_3_21;
wire din_valid_3_21;
wire [63:0] din_3_22;
wire din_valid_3_22;
wire [63:0] din_3_23;
wire din_valid_3_23;
wire [63:0] din_3_24;
wire din_valid_3_24;
wire [63:0] din_3_25;
wire din_valid_3_25;
wire [63:0] din_3_26;
wire din_valid_3_26;
wire [63:0] din_3_27;
wire din_valid_3_27;
wire [63:0] din_3_28;
wire din_valid_3_28;
wire [63:0] din_3_29;
wire din_valid_3_29;
wire [63:0] din_3_30;
wire din_valid_3_30;
wire [63:0] din_3_31;
wire din_valid_3_31;
wire [63:0] din_4_0;
wire din_valid_4_0;
wire [63:0] din_4_1;
wire din_valid_4_1;
wire [63:0] din_4_2;
wire din_valid_4_2;
wire [63:0] din_4_3;
wire din_valid_4_3;
wire [63:0] din_4_4;
wire din_valid_4_4;
wire [63:0] din_4_5;
wire din_valid_4_5;
wire [63:0] din_4_6;
wire din_valid_4_6;
wire [63:0] din_4_7;
wire din_valid_4_7;
wire [63:0] din_4_8;
wire din_valid_4_8;
wire [63:0] din_4_9;
wire din_valid_4_9;
wire [63:0] din_4_10;
wire din_valid_4_10;
wire [63:0] din_4_11;
wire din_valid_4_11;
wire [63:0] din_4_12;
wire din_valid_4_12;
wire [63:0] din_4_13;
wire din_valid_4_13;
wire [63:0] din_4_14;
wire din_valid_4_14;
wire [63:0] din_4_15;
wire din_valid_4_15;
wire [63:0] din_4_16;
wire din_valid_4_16;
wire [63:0] din_4_17;
wire din_valid_4_17;
wire [63:0] din_4_18;
wire din_valid_4_18;
wire [63:0] din_4_19;
wire din_valid_4_19;
wire [63:0] din_4_20;
wire din_valid_4_20;
wire [63:0] din_4_21;
wire din_valid_4_21;
wire [63:0] din_4_22;
wire din_valid_4_22;
wire [63:0] din_4_23;
wire din_valid_4_23;
wire [63:0] din_4_24;
wire din_valid_4_24;
wire [63:0] din_4_25;
wire din_valid_4_25;
wire [63:0] din_4_26;
wire din_valid_4_26;
wire [63:0] din_4_27;
wire din_valid_4_27;
wire [63:0] din_4_28;
wire din_valid_4_28;
wire [63:0] din_4_29;
wire din_valid_4_29;
wire [63:0] din_4_30;
wire din_valid_4_30;
wire [63:0] din_4_31;
wire din_valid_4_31;
wire [63:0] din_5_0;
wire din_valid_5_0;
wire [63:0] din_5_1;
wire din_valid_5_1;
wire [63:0] din_5_2;
wire din_valid_5_2;
wire [63:0] din_5_3;
wire din_valid_5_3;
wire [63:0] din_5_4;
wire din_valid_5_4;
wire [63:0] din_5_5;
wire din_valid_5_5;
wire [63:0] din_5_6;
wire din_valid_5_6;
wire [63:0] din_5_7;
wire din_valid_5_7;
wire [63:0] din_5_8;
wire din_valid_5_8;
wire [63:0] din_5_9;
wire din_valid_5_9;
wire [63:0] din_5_10;
wire din_valid_5_10;
wire [63:0] din_5_11;
wire din_valid_5_11;
wire [63:0] din_5_12;
wire din_valid_5_12;
wire [63:0] din_5_13;
wire din_valid_5_13;
wire [63:0] din_5_14;
wire din_valid_5_14;
wire [63:0] din_5_15;
wire din_valid_5_15;
wire [63:0] din_5_16;
wire din_valid_5_16;
wire [63:0] din_5_17;
wire din_valid_5_17;
wire [63:0] din_5_18;
wire din_valid_5_18;
wire [63:0] din_5_19;
wire din_valid_5_19;
wire [63:0] din_5_20;
wire din_valid_5_20;
wire [63:0] din_5_21;
wire din_valid_5_21;
wire [63:0] din_5_22;
wire din_valid_5_22;
wire [63:0] din_5_23;
wire din_valid_5_23;
wire [63:0] din_5_24;
wire din_valid_5_24;
wire [63:0] din_5_25;
wire din_valid_5_25;
wire [63:0] din_5_26;
wire din_valid_5_26;
wire [63:0] din_5_27;
wire din_valid_5_27;
wire [63:0] din_5_28;
wire din_valid_5_28;
wire [63:0] din_5_29;
wire din_valid_5_29;
wire [63:0] din_5_30;
wire din_valid_5_30;
wire [63:0] din_5_31;
wire din_valid_5_31;
wire [63:0] din_6_0;
wire din_valid_6_0;
wire [63:0] din_6_1;
wire din_valid_6_1;
wire [63:0] din_6_2;
wire din_valid_6_2;
wire [63:0] din_6_3;
wire din_valid_6_3;
wire [63:0] din_6_4;
wire din_valid_6_4;
wire [63:0] din_6_5;
wire din_valid_6_5;
wire [63:0] din_6_6;
wire din_valid_6_6;
wire [63:0] din_6_7;
wire din_valid_6_7;
wire [63:0] din_6_8;
wire din_valid_6_8;
wire [63:0] din_6_9;
wire din_valid_6_9;
wire [63:0] din_6_10;
wire din_valid_6_10;
wire [63:0] din_6_11;
wire din_valid_6_11;
wire [63:0] din_6_12;
wire din_valid_6_12;
wire [63:0] din_6_13;
wire din_valid_6_13;
wire [63:0] din_6_14;
wire din_valid_6_14;
wire [63:0] din_6_15;
wire din_valid_6_15;
wire [63:0] din_6_16;
wire din_valid_6_16;
wire [63:0] din_6_17;
wire din_valid_6_17;
wire [63:0] din_6_18;
wire din_valid_6_18;
wire [63:0] din_6_19;
wire din_valid_6_19;
wire [63:0] din_6_20;
wire din_valid_6_20;
wire [63:0] din_6_21;
wire din_valid_6_21;
wire [63:0] din_6_22;
wire din_valid_6_22;
wire [63:0] din_6_23;
wire din_valid_6_23;
wire [63:0] din_6_24;
wire din_valid_6_24;
wire [63:0] din_6_25;
wire din_valid_6_25;
wire [63:0] din_6_26;
wire din_valid_6_26;
wire [63:0] din_6_27;
wire din_valid_6_27;
wire [63:0] din_6_28;
wire din_valid_6_28;
wire [63:0] din_6_29;
wire din_valid_6_29;
wire [63:0] din_6_30;
wire din_valid_6_30;
wire [63:0] din_6_31;
wire din_valid_6_31;
wire [63:0] din_7_0;
wire din_valid_7_0;
wire [63:0] din_7_1;
wire din_valid_7_1;
wire [63:0] din_7_2;
wire din_valid_7_2;
wire [63:0] din_7_3;
wire din_valid_7_3;
wire [63:0] din_7_4;
wire din_valid_7_4;
wire [63:0] din_7_5;
wire din_valid_7_5;
wire [63:0] din_7_6;
wire din_valid_7_6;
wire [63:0] din_7_7;
wire din_valid_7_7;
wire [63:0] din_7_8;
wire din_valid_7_8;
wire [63:0] din_7_9;
wire din_valid_7_9;
wire [63:0] din_7_10;
wire din_valid_7_10;
wire [63:0] din_7_11;
wire din_valid_7_11;
wire [63:0] din_7_12;
wire din_valid_7_12;
wire [63:0] din_7_13;
wire din_valid_7_13;
wire [63:0] din_7_14;
wire din_valid_7_14;
wire [63:0] din_7_15;
wire din_valid_7_15;
wire [63:0] din_7_16;
wire din_valid_7_16;
wire [63:0] din_7_17;
wire din_valid_7_17;
wire [63:0] din_7_18;
wire din_valid_7_18;
wire [63:0] din_7_19;
wire din_valid_7_19;
wire [63:0] din_7_20;
wire din_valid_7_20;
wire [63:0] din_7_21;
wire din_valid_7_21;
wire [63:0] din_7_22;
wire din_valid_7_22;
wire [63:0] din_7_23;
wire din_valid_7_23;
wire [63:0] din_7_24;
wire din_valid_7_24;
wire [63:0] din_7_25;
wire din_valid_7_25;
wire [63:0] din_7_26;
wire din_valid_7_26;
wire [63:0] din_7_27;
wire din_valid_7_27;
wire [63:0] din_7_28;
wire din_valid_7_28;
wire [63:0] din_7_29;
wire din_valid_7_29;
wire [63:0] din_7_30;
wire din_valid_7_30;
wire [63:0] din_7_31;
wire din_valid_7_31;

reg [63:0] din_reg;
reg din_valid_reg;

assign din_0_0 = {din[7:0],din_reg[63:8]};
assign din_0_1 = {din[15:0],din_reg[63:16]};
assign din_0_2 = {din[23:0],din_reg[63:24]};
assign din_0_3 = {din[31:0],din_reg[63:32]};
assign din_0_4 = {din[39:0],din_reg[63:40]};
assign din_0_5 = {din[47:0],din_reg[63:48]};
assign din_0_6 = {din[55:0],din_reg[63:56]};

assign din_0_7 = din[63:0];
assign din_0_8 = din[71:8];
assign din_0_9 = din[79:16];
assign din_0_10 = din[87:24];
assign din_0_11 = din[95:32];
assign din_0_12 = din[103:40];
assign din_0_13 = din[111:48];
assign din_0_14 = din[119:56];
assign din_0_15 = din[127:64];
assign din_0_16 = din[135:72];
assign din_0_17 = din[143:80];
assign din_0_18 = din[151:88];
assign din_0_19 = din[159:96];
assign din_0_20 = din[167:104];
assign din_0_21 = din[175:112];
assign din_0_22 = din[183:120];
assign din_0_23 = din[191:128];
assign din_0_24 = din[199:136];
assign din_0_25 = din[207:144];
assign din_0_26 = din[215:152];
assign din_0_27 = din[223:160];
assign din_0_28 = din[231:168];
assign din_0_29 = din[239:176];
assign din_0_30 = din[247:184];
assign din_0_31 = din[255:192];
assign din_1_0 = {din[7:0],din_reg[63:8]};
assign din_1_1 = {din[15:0],din_reg[63:16]};
assign din_1_2 = {din[23:0],din_reg[63:24]};
assign din_1_3 = {din[31:0],din_reg[63:32]};
assign din_1_4 = {din[39:0],din_reg[63:40]};
assign din_1_5 = {din[47:0],din_reg[63:48]};
assign din_1_6 = {din[55:0],din_reg[63:56]};

assign din_1_7 = din[63:0];
assign din_1_8 = din[71:8];
assign din_1_9 = din[79:16];
assign din_1_10 = din[87:24];
assign din_1_11 = din[95:32];
assign din_1_12 = din[103:40];
assign din_1_13 = din[111:48];
assign din_1_14 = din[119:56];
assign din_1_15 = din[127:64];
assign din_1_16 = din[135:72];
assign din_1_17 = din[143:80];
assign din_1_18 = din[151:88];
assign din_1_19 = din[159:96];
assign din_1_20 = din[167:104];
assign din_1_21 = din[175:112];
assign din_1_22 = din[183:120];
assign din_1_23 = din[191:128];
assign din_1_24 = din[199:136];
assign din_1_25 = din[207:144];
assign din_1_26 = din[215:152];
assign din_1_27 = din[223:160];
assign din_1_28 = din[231:168];
assign din_1_29 = din[239:176];
assign din_1_30 = din[247:184];
assign din_1_31 = din[255:192];
assign din_2_0 = {din[7:0],din_reg[63:8]};
assign din_2_1 = {din[15:0],din_reg[63:16]};
assign din_2_2 = {din[23:0],din_reg[63:24]};
assign din_2_3 = {din[31:0],din_reg[63:32]};
assign din_2_4 = {din[39:0],din_reg[63:40]};
assign din_2_5 = {din[47:0],din_reg[63:48]};
assign din_2_6 = {din[55:0],din_reg[63:56]};

assign din_2_7 = din[63:0];
assign din_2_8 = din[71:8];
assign din_2_9 = din[79:16];
assign din_2_10 = din[87:24];
assign din_2_11 = din[95:32];
assign din_2_12 = din[103:40];
assign din_2_13 = din[111:48];
assign din_2_14 = din[119:56];
assign din_2_15 = din[127:64];
assign din_2_16 = din[135:72];
assign din_2_17 = din[143:80];
assign din_2_18 = din[151:88];
assign din_2_19 = din[159:96];
assign din_2_20 = din[167:104];
assign din_2_21 = din[175:112];
assign din_2_22 = din[183:120];
assign din_2_23 = din[191:128];
assign din_2_24 = din[199:136];
assign din_2_25 = din[207:144];
assign din_2_26 = din[215:152];
assign din_2_27 = din[223:160];
assign din_2_28 = din[231:168];
assign din_2_29 = din[239:176];
assign din_2_30 = din[247:184];
assign din_2_31 = din[255:192];
assign din_3_0 = {din[7:0],din_reg[63:8]};
assign din_3_1 = {din[15:0],din_reg[63:16]};
assign din_3_2 = {din[23:0],din_reg[63:24]};
assign din_3_3 = {din[31:0],din_reg[63:32]};
assign din_3_4 = {din[39:0],din_reg[63:40]};
assign din_3_5 = {din[47:0],din_reg[63:48]};
assign din_3_6 = {din[55:0],din_reg[63:56]};

assign din_3_7 = din[63:0];
assign din_3_8 = din[71:8];
assign din_3_9 = din[79:16];
assign din_3_10 = din[87:24];
assign din_3_11 = din[95:32];
assign din_3_12 = din[103:40];
assign din_3_13 = din[111:48];
assign din_3_14 = din[119:56];
assign din_3_15 = din[127:64];
assign din_3_16 = din[135:72];
assign din_3_17 = din[143:80];
assign din_3_18 = din[151:88];
assign din_3_19 = din[159:96];
assign din_3_20 = din[167:104];
assign din_3_21 = din[175:112];
assign din_3_22 = din[183:120];
assign din_3_23 = din[191:128];
assign din_3_24 = din[199:136];
assign din_3_25 = din[207:144];
assign din_3_26 = din[215:152];
assign din_3_27 = din[223:160];
assign din_3_28 = din[231:168];
assign din_3_29 = din[239:176];
assign din_3_30 = din[247:184];
assign din_3_31 = din[255:192];
assign din_4_0 = {din[7:0],din_reg[63:8]};
assign din_4_1 = {din[15:0],din_reg[63:16]};
assign din_4_2 = {din[23:0],din_reg[63:24]};
assign din_4_3 = {din[31:0],din_reg[63:32]};
assign din_4_4 = {din[39:0],din_reg[63:40]};
assign din_4_5 = {din[47:0],din_reg[63:48]};
assign din_4_6 = {din[55:0],din_reg[63:56]};

assign din_4_7 = din[63:0];
assign din_4_8 = din[71:8];
assign din_4_9 = din[79:16];
assign din_4_10 = din[87:24];
assign din_4_11 = din[95:32];
assign din_4_12 = din[103:40];
assign din_4_13 = din[111:48];
assign din_4_14 = din[119:56];
assign din_4_15 = din[127:64];
assign din_4_16 = din[135:72];
assign din_4_17 = din[143:80];
assign din_4_18 = din[151:88];
assign din_4_19 = din[159:96];
assign din_4_20 = din[167:104];
assign din_4_21 = din[175:112];
assign din_4_22 = din[183:120];
assign din_4_23 = din[191:128];
assign din_4_24 = din[199:136];
assign din_4_25 = din[207:144];
assign din_4_26 = din[215:152];
assign din_4_27 = din[223:160];
assign din_4_28 = din[231:168];
assign din_4_29 = din[239:176];
assign din_4_30 = din[247:184];
assign din_4_31 = din[255:192];
assign din_5_0 = {din[7:0],din_reg[63:8]};
assign din_5_1 = {din[15:0],din_reg[63:16]};
assign din_5_2 = {din[23:0],din_reg[63:24]};
assign din_5_3 = {din[31:0],din_reg[63:32]};
assign din_5_4 = {din[39:0],din_reg[63:40]};
assign din_5_5 = {din[47:0],din_reg[63:48]};
assign din_5_6 = {din[55:0],din_reg[63:56]};

assign din_5_7 = din[63:0];
assign din_5_8 = din[71:8];
assign din_5_9 = din[79:16];
assign din_5_10 = din[87:24];
assign din_5_11 = din[95:32];
assign din_5_12 = din[103:40];
assign din_5_13 = din[111:48];
assign din_5_14 = din[119:56];
assign din_5_15 = din[127:64];
assign din_5_16 = din[135:72];
assign din_5_17 = din[143:80];
assign din_5_18 = din[151:88];
assign din_5_19 = din[159:96];
assign din_5_20 = din[167:104];
assign din_5_21 = din[175:112];
assign din_5_22 = din[183:120];
assign din_5_23 = din[191:128];
assign din_5_24 = din[199:136];
assign din_5_25 = din[207:144];
assign din_5_26 = din[215:152];
assign din_5_27 = din[223:160];
assign din_5_28 = din[231:168];
assign din_5_29 = din[239:176];
assign din_5_30 = din[247:184];
assign din_5_31 = din[255:192];
assign din_6_0 = {din[7:0],din_reg[63:8]};
assign din_6_1 = {din[15:0],din_reg[63:16]};
assign din_6_2 = {din[23:0],din_reg[63:24]};
assign din_6_3 = {din[31:0],din_reg[63:32]};
assign din_6_4 = {din[39:0],din_reg[63:40]};
assign din_6_5 = {din[47:0],din_reg[63:48]};
assign din_6_6 = {din[55:0],din_reg[63:56]};

assign din_6_7 = din[63:0];
assign din_6_8 = din[71:8];
assign din_6_9 = din[79:16];
assign din_6_10 = din[87:24];
assign din_6_11 = din[95:32];
assign din_6_12 = din[103:40];
assign din_6_13 = din[111:48];
assign din_6_14 = din[119:56];
assign din_6_15 = din[127:64];
assign din_6_16 = din[135:72];
assign din_6_17 = din[143:80];
assign din_6_18 = din[151:88];
assign din_6_19 = din[159:96];
assign din_6_20 = din[167:104];
assign din_6_21 = din[175:112];
assign din_6_22 = din[183:120];
assign din_6_23 = din[191:128];
assign din_6_24 = din[199:136];
assign din_6_25 = din[207:144];
assign din_6_26 = din[215:152];
assign din_6_27 = din[223:160];
assign din_6_28 = din[231:168];
assign din_6_29 = din[239:176];
assign din_6_30 = din[247:184];
assign din_6_31 = din[255:192];
assign din_7_0 = {din[7:0],din_reg[63:8]};
assign din_7_1 = {din[15:0],din_reg[63:16]};
assign din_7_2 = {din[23:0],din_reg[63:24]};
assign din_7_3 = {din[31:0],din_reg[63:32]};
assign din_7_4 = {din[39:0],din_reg[63:40]};
assign din_7_5 = {din[47:0],din_reg[63:48]};
assign din_7_6 = {din[55:0],din_reg[63:56]};

assign din_7_7 = din[63:0];
assign din_7_8 = din[71:8];
assign din_7_9 = din[79:16];
assign din_7_10 = din[87:24];
assign din_7_11 = din[95:32];
assign din_7_12 = din[103:40];
assign din_7_13 = din[111:48];
assign din_7_14 = din[119:56];
assign din_7_15 = din[127:64];
assign din_7_16 = din[135:72];
assign din_7_17 = din[143:80];
assign din_7_18 = din[151:88];
assign din_7_19 = din[159:96];
assign din_7_20 = din[167:104];
assign din_7_21 = din[175:112];
assign din_7_22 = din[183:120];
assign din_7_23 = din[191:128];
assign din_7_24 = din[199:136];
assign din_7_25 = din[207:144];
assign din_7_26 = din[215:152];
assign din_7_27 = din[223:160];
assign din_7_28 = din[231:168];
assign din_7_29 = din[239:176];
assign din_7_30 = din[247:184];
assign din_7_31 = din[255:192];

//Valid signals
assign din_valid_0_0 = din_valid & din_valid_reg;
assign din_valid_1_0 = din_valid & din_valid_reg;
assign din_valid_0_1 = din_valid & din_valid_reg;
assign din_valid_1_1 = din_valid & din_valid_reg;
assign din_valid_0_2 = din_valid & din_valid_reg;
assign din_valid_1_2 = din_valid & din_valid_reg;
assign din_valid_0_3 = din_valid & din_valid_reg;
assign din_valid_1_3 = din_valid & din_valid_reg;
assign din_valid_0_4 = din_valid & din_valid_reg;
assign din_valid_1_4 = din_valid & din_valid_reg;
assign din_valid_0_5 = din_valid & din_valid_reg;
assign din_valid_1_5 = din_valid & din_valid_reg;
assign din_valid_0_6 = din_valid & din_valid_reg;
assign din_valid_1_6 = din_valid & din_valid_reg;
assign din_valid_0_7 = din_valid;
assign din_valid_1_7 = din_valid;
assign din_valid_0_8 = din_valid;
assign din_valid_1_8 = din_valid;
assign din_valid_0_9 = din_valid;
assign din_valid_1_9 = din_valid;
assign din_valid_0_10 = din_valid;
assign din_valid_1_10 = din_valid;
assign din_valid_0_11 = din_valid;
assign din_valid_1_11 = din_valid;
assign din_valid_0_12 = din_valid;
assign din_valid_1_12 = din_valid;
assign din_valid_0_13 = din_valid;
assign din_valid_1_13 = din_valid;
assign din_valid_0_14 = din_valid;
assign din_valid_1_14 = din_valid;
assign din_valid_0_15 = din_valid;
assign din_valid_1_15 = din_valid;
assign din_valid_0_16 = din_valid;
assign din_valid_1_16 = din_valid;
assign din_valid_0_17 = din_valid;
assign din_valid_1_17 = din_valid;
assign din_valid_0_18 = din_valid;
assign din_valid_1_18 = din_valid;
assign din_valid_0_19 = din_valid;
assign din_valid_1_19 = din_valid;
assign din_valid_0_20 = din_valid;
assign din_valid_1_20 = din_valid;
assign din_valid_0_21 = din_valid;
assign din_valid_1_21 = din_valid;
assign din_valid_0_22 = din_valid;
assign din_valid_1_22 = din_valid;
assign din_valid_0_23 = din_valid;
assign din_valid_1_23 = din_valid;
assign din_valid_0_24 = din_valid;
assign din_valid_1_24 = din_valid;
assign din_valid_0_25 = din_valid;
assign din_valid_1_25 = din_valid;
assign din_valid_0_26 = din_valid;
assign din_valid_1_26 = din_valid;
assign din_valid_0_27 = din_valid;
assign din_valid_1_27 = din_valid;
assign din_valid_0_28 = din_valid;
assign din_valid_1_28 = din_valid;
assign din_valid_0_29 = din_valid;
assign din_valid_1_29 = din_valid;
assign din_valid_0_30 = din_valid;
assign din_valid_1_30 = din_valid;
assign din_valid_0_31 = din_valid;
assign din_valid_1_31 = din_valid;

assign din_valid_2_0 = din_valid & din_valid_reg;
assign din_valid_2_1 = din_valid & din_valid_reg;
assign din_valid_2_2 = din_valid & din_valid_reg;
assign din_valid_2_3 = din_valid & din_valid_reg;
assign din_valid_2_4 = din_valid & din_valid_reg;
assign din_valid_2_5 = din_valid & din_valid_reg;
assign din_valid_2_6 = din_valid;
assign din_valid_2_7 = din_valid;
assign din_valid_2_8 = din_valid;
assign din_valid_2_9 = din_valid;
assign din_valid_2_10 = din_valid;
assign din_valid_2_11 = din_valid;
assign din_valid_2_12 = din_valid;
assign din_valid_2_13 = din_valid;
assign din_valid_2_14 = din_valid;
assign din_valid_2_15 = din_valid;
assign din_valid_2_16 = din_valid;
assign din_valid_2_17 = din_valid;
assign din_valid_2_18 = din_valid;
assign din_valid_2_19 = din_valid;
assign din_valid_2_20 = din_valid;
assign din_valid_2_21 = din_valid;
assign din_valid_2_22 = din_valid;
assign din_valid_2_23 = din_valid;
assign din_valid_2_24 = din_valid;
assign din_valid_2_25 = din_valid;
assign din_valid_2_26 = din_valid;
assign din_valid_2_27 = din_valid;
assign din_valid_2_28 = din_valid;
assign din_valid_2_29 = din_valid;
assign din_valid_2_30 = din_valid;
assign din_valid_2_31 = din_valid;

assign din_valid_3_0 = din_valid & din_valid_reg;
assign din_valid_3_1 = din_valid & din_valid_reg;
assign din_valid_3_2 = din_valid & din_valid_reg;
assign din_valid_3_3 = din_valid & din_valid_reg;
assign din_valid_3_4 = din_valid & din_valid_reg;
assign din_valid_3_5 = din_valid;
assign din_valid_3_6 = din_valid;
assign din_valid_3_7 = din_valid;
assign din_valid_3_8 = din_valid;
assign din_valid_3_9 = din_valid;
assign din_valid_3_10 = din_valid;
assign din_valid_3_11 = din_valid;
assign din_valid_3_12 = din_valid;
assign din_valid_3_13 = din_valid;
assign din_valid_3_14 = din_valid;
assign din_valid_3_15 = din_valid;
assign din_valid_3_16 = din_valid;
assign din_valid_3_17 = din_valid;
assign din_valid_3_18 = din_valid;
assign din_valid_3_19 = din_valid;
assign din_valid_3_20 = din_valid;
assign din_valid_3_21 = din_valid;
assign din_valid_3_22 = din_valid;
assign din_valid_3_23 = din_valid;
assign din_valid_3_24 = din_valid;
assign din_valid_3_25 = din_valid;
assign din_valid_3_26 = din_valid;
assign din_valid_3_27 = din_valid;
assign din_valid_3_28 = din_valid;
assign din_valid_3_29 = din_valid;
assign din_valid_3_30 = din_valid;
assign din_valid_3_31 = din_valid;

assign din_valid_4_0 = din_valid & din_valid_reg;
assign din_valid_4_1 = din_valid & din_valid_reg;
assign din_valid_4_2 = din_valid & din_valid_reg;
assign din_valid_4_3 = din_valid & din_valid_reg;
assign din_valid_4_4 = din_valid;
assign din_valid_4_5 = din_valid;
assign din_valid_4_6 = din_valid;
assign din_valid_4_7 = din_valid;
assign din_valid_4_8 = din_valid;
assign din_valid_4_9 = din_valid;
assign din_valid_4_10 = din_valid;
assign din_valid_4_11 = din_valid;
assign din_valid_4_12 = din_valid;
assign din_valid_4_13 = din_valid;
assign din_valid_4_14 = din_valid;
assign din_valid_4_15 = din_valid;
assign din_valid_4_16 = din_valid;
assign din_valid_4_17 = din_valid;
assign din_valid_4_18 = din_valid;
assign din_valid_4_19 = din_valid;
assign din_valid_4_20 = din_valid;
assign din_valid_4_21 = din_valid;
assign din_valid_4_22 = din_valid;
assign din_valid_4_23 = din_valid;
assign din_valid_4_24 = din_valid;
assign din_valid_4_25 = din_valid;
assign din_valid_4_26 = din_valid;
assign din_valid_4_27 = din_valid;
assign din_valid_4_28 = din_valid;
assign din_valid_4_29 = din_valid;
assign din_valid_4_30 = din_valid;
assign din_valid_4_31 = din_valid;

assign din_valid_5_0 = din_valid & din_valid_reg;
assign din_valid_5_1 = din_valid & din_valid_reg;
assign din_valid_5_2 = din_valid & din_valid_reg;
assign din_valid_5_3 = din_valid;
assign din_valid_5_4 = din_valid;
assign din_valid_5_5 = din_valid;
assign din_valid_5_6 = din_valid;
assign din_valid_5_7 = din_valid;
assign din_valid_5_8 = din_valid;
assign din_valid_5_9 = din_valid;
assign din_valid_5_10 = din_valid;
assign din_valid_5_11 = din_valid;
assign din_valid_5_12 = din_valid;
assign din_valid_5_13 = din_valid;
assign din_valid_5_14 = din_valid;
assign din_valid_5_15 = din_valid;
assign din_valid_5_16 = din_valid;
assign din_valid_5_17 = din_valid;
assign din_valid_5_18 = din_valid;
assign din_valid_5_19 = din_valid;
assign din_valid_5_20 = din_valid;
assign din_valid_5_21 = din_valid;
assign din_valid_5_22 = din_valid;
assign din_valid_5_23 = din_valid;
assign din_valid_5_24 = din_valid;
assign din_valid_5_25 = din_valid;
assign din_valid_5_26 = din_valid;
assign din_valid_5_27 = din_valid;
assign din_valid_5_28 = din_valid;
assign din_valid_5_29 = din_valid;
assign din_valid_5_30 = din_valid;
assign din_valid_5_31 = din_valid;

assign din_valid_6_0 = din_valid & din_valid_reg;
assign din_valid_6_1 = din_valid & din_valid_reg;
assign din_valid_6_2 = din_valid;
assign din_valid_6_3 = din_valid;
assign din_valid_6_4 = din_valid;
assign din_valid_6_5 = din_valid;
assign din_valid_6_6 = din_valid;
assign din_valid_6_7 = din_valid;
assign din_valid_6_8 = din_valid;
assign din_valid_6_9 = din_valid;
assign din_valid_6_10 = din_valid;
assign din_valid_6_11 = din_valid;
assign din_valid_6_12 = din_valid;
assign din_valid_6_13 = din_valid;
assign din_valid_6_14 = din_valid;
assign din_valid_6_15 = din_valid;
assign din_valid_6_16 = din_valid;
assign din_valid_6_17 = din_valid;
assign din_valid_6_18 = din_valid;
assign din_valid_6_19 = din_valid;
assign din_valid_6_20 = din_valid;
assign din_valid_6_21 = din_valid;
assign din_valid_6_22 = din_valid;
assign din_valid_6_23 = din_valid;
assign din_valid_6_24 = din_valid;
assign din_valid_6_25 = din_valid;
assign din_valid_6_26 = din_valid;
assign din_valid_6_27 = din_valid;
assign din_valid_6_28 = din_valid;
assign din_valid_6_29 = din_valid;
assign din_valid_6_30 = din_valid;
assign din_valid_6_31 = din_valid;

assign din_valid_7_0 = din_valid & din_valid_reg;
assign din_valid_7_1 = din_valid;
assign din_valid_7_2 = din_valid;
assign din_valid_7_3 = din_valid;
assign din_valid_7_4 = din_valid;
assign din_valid_7_5 = din_valid;
assign din_valid_7_6 = din_valid;
assign din_valid_7_7 = din_valid;
assign din_valid_7_8 = din_valid;
assign din_valid_7_9 = din_valid;
assign din_valid_7_10 = din_valid;
assign din_valid_7_11 = din_valid;
assign din_valid_7_12 = din_valid;
assign din_valid_7_13 = din_valid;
assign din_valid_7_14 = din_valid;
assign din_valid_7_15 = din_valid;
assign din_valid_7_16 = din_valid;
assign din_valid_7_17 = din_valid;
assign din_valid_7_18 = din_valid;
assign din_valid_7_19 = din_valid;
assign din_valid_7_20 = din_valid;
assign din_valid_7_21 = din_valid;
assign din_valid_7_22 = din_valid;
assign din_valid_7_23 = din_valid;
assign din_valid_7_24 = din_valid;
assign din_valid_7_25 = din_valid;
assign din_valid_7_26 = din_valid;
assign din_valid_7_27 = din_valid;
assign din_valid_7_28 = din_valid;
assign din_valid_7_29 = din_valid;
assign din_valid_7_30 = din_valid;
assign din_valid_7_31 = din_valid;


always @ (posedge clk) begin
    //din_reg <= din[127:64];
    din_reg <= din[255:192];
    din_valid_reg <= din_valid;
end


hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_0 (
	.clk (clk),
	.din0 (din_0_0),
	.din0_valid (din_valid_0_0),
	.din1 (din_0_1),
	.din1_valid (din_valid_0_1),
	.dout0 (dout_0_0),
	.dout0_valid (dout_valid_0_0),
	.dout1 (dout_0_1),
	.dout1_valid (dout_valid_0_1)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_1 (
	.clk (clk),
	.din0 (din_0_2),
	.din0_valid (din_valid_0_2),
	.din1 (din_0_3),
	.din1_valid (din_valid_0_3),
	.dout0 (dout_0_2),
	.dout0_valid (dout_valid_0_2),
	.dout1 (dout_0_3),
	.dout1_valid (dout_valid_0_3)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_2 (
	.clk (clk),
	.din0 (din_0_4),
	.din0_valid (din_valid_0_4),
	.din1 (din_0_5),
	.din1_valid (din_valid_0_5),
	.dout0 (dout_0_4),
	.dout0_valid (dout_valid_0_4),
	.dout1 (dout_0_5),
	.dout1_valid (dout_valid_0_5)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_3 (
	.clk (clk),
	.din0 (din_0_6),
	.din0_valid (din_valid_0_6),
	.din1 (din_0_7),
	.din1_valid (din_valid_0_7),
	.dout0 (dout_0_6),
	.dout0_valid (dout_valid_0_6),
	.dout1 (dout_0_7),
	.dout1_valid (dout_valid_0_7)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_4 (
	.clk (clk),
	.din0 (din_0_8),
	.din0_valid (din_valid_0_8),
	.din1 (din_0_9),
	.din1_valid (din_valid_0_9),
	.dout0 (dout_0_8),
	.dout0_valid (dout_valid_0_8),
	.dout1 (dout_0_9),
	.dout1_valid (dout_valid_0_9)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_5 (
	.clk (clk),
	.din0 (din_0_10),
	.din0_valid (din_valid_0_10),
	.din1 (din_0_11),
	.din1_valid (din_valid_0_11),
	.dout0 (dout_0_10),
	.dout0_valid (dout_valid_0_10),
	.dout1 (dout_0_11),
	.dout1_valid (dout_valid_0_11)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_6 (
	.clk (clk),
	.din0 (din_0_12),
	.din0_valid (din_valid_0_12),
	.din1 (din_0_13),
	.din1_valid (din_valid_0_13),
	.dout0 (dout_0_12),
	.dout0_valid (dout_valid_0_12),
	.dout1 (dout_0_13),
	.dout1_valid (dout_valid_0_13)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_7 (
	.clk (clk),
	.din0 (din_0_14),
	.din0_valid (din_valid_0_14),
	.din1 (din_0_15),
	.din1_valid (din_valid_0_15),
	.dout0 (dout_0_14),
	.dout0_valid (dout_valid_0_14),
	.dout1 (dout_0_15),
	.dout1_valid (dout_valid_0_15)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_8 (
	.clk (clk),
	.din0 (din_0_16),
	.din0_valid (din_valid_0_16),
	.din1 (din_0_17),
	.din1_valid (din_valid_0_17),
	.dout0 (dout_0_16),
	.dout0_valid (dout_valid_0_16),
	.dout1 (dout_0_17),
	.dout1_valid (dout_valid_0_17)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_9 (
	.clk (clk),
	.din0 (din_0_18),
	.din0_valid (din_valid_0_18),
	.din1 (din_0_19),
	.din1_valid (din_valid_0_19),
	.dout0 (dout_0_18),
	.dout0_valid (dout_valid_0_18),
	.dout1 (dout_0_19),
	.dout1_valid (dout_valid_0_19)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_10 (
	.clk (clk),
	.din0 (din_0_20),
	.din0_valid (din_valid_0_20),
	.din1 (din_0_21),
	.din1_valid (din_valid_0_21),
	.dout0 (dout_0_20),
	.dout0_valid (dout_valid_0_20),
	.dout1 (dout_0_21),
	.dout1_valid (dout_valid_0_21)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_11 (
	.clk (clk),
	.din0 (din_0_22),
	.din0_valid (din_valid_0_22),
	.din1 (din_0_23),
	.din1_valid (din_valid_0_23),
	.dout0 (dout_0_22),
	.dout0_valid (dout_valid_0_22),
	.dout1 (dout_0_23),
	.dout1_valid (dout_valid_0_23)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_12 (
	.clk (clk),
	.din0 (din_0_24),
	.din0_valid (din_valid_0_24),
	.din1 (din_0_25),
	.din1_valid (din_valid_0_25),
	.dout0 (dout_0_24),
	.dout0_valid (dout_valid_0_24),
	.dout1 (dout_0_25),
	.dout1_valid (dout_valid_0_25)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_13 (
	.clk (clk),
	.din0 (din_0_26),
	.din0_valid (din_valid_0_26),
	.din1 (din_0_27),
	.din1_valid (din_valid_0_27),
	.dout0 (dout_0_26),
	.dout0_valid (dout_valid_0_26),
	.dout1 (dout_0_27),
	.dout1_valid (dout_valid_0_27)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_14 (
	.clk (clk),
	.din0 (din_0_28),
	.din0_valid (din_valid_0_28),
	.din1 (din_0_29),
	.din1_valid (din_valid_0_29),
	.dout0 (dout_0_28),
	.dout0_valid (dout_valid_0_28),
	.dout1 (dout_0_29),
	.dout1_valid (dout_valid_0_29)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap0.mif")
)
hashtable_0_15 (
	.clk (clk),
	.din0 (din_0_30),
	.din0_valid (din_valid_0_30),
	.din1 (din_0_31),
	.din1_valid (din_valid_0_31),
	.dout0 (dout_0_30),
	.dout0_valid (dout_valid_0_30),
	.dout1 (dout_0_31),
	.dout1_valid (dout_valid_0_31)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_0 (
	.clk (clk),
	.din0 (din_1_0),
	.din0_valid (din_valid_1_0),
	.din1 (din_1_1),
	.din1_valid (din_valid_1_1),
	.dout0 (dout_1_0),
	.dout0_valid (dout_valid_1_0),
	.dout1 (dout_1_1),
	.dout1_valid (dout_valid_1_1)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_1 (
	.clk (clk),
	.din0 (din_1_2),
	.din0_valid (din_valid_1_2),
	.din1 (din_1_3),
	.din1_valid (din_valid_1_3),
	.dout0 (dout_1_2),
	.dout0_valid (dout_valid_1_2),
	.dout1 (dout_1_3),
	.dout1_valid (dout_valid_1_3)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_2 (
	.clk (clk),
	.din0 (din_1_4),
	.din0_valid (din_valid_1_4),
	.din1 (din_1_5),
	.din1_valid (din_valid_1_5),
	.dout0 (dout_1_4),
	.dout0_valid (dout_valid_1_4),
	.dout1 (dout_1_5),
	.dout1_valid (dout_valid_1_5)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_3 (
	.clk (clk),
	.din0 (din_1_6),
	.din0_valid (din_valid_1_6),
	.din1 (din_1_7),
	.din1_valid (din_valid_1_7),
	.dout0 (dout_1_6),
	.dout0_valid (dout_valid_1_6),
	.dout1 (dout_1_7),
	.dout1_valid (dout_valid_1_7)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_4 (
	.clk (clk),
	.din0 (din_1_8),
	.din0_valid (din_valid_1_8),
	.din1 (din_1_9),
	.din1_valid (din_valid_1_9),
	.dout0 (dout_1_8),
	.dout0_valid (dout_valid_1_8),
	.dout1 (dout_1_9),
	.dout1_valid (dout_valid_1_9)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_5 (
	.clk (clk),
	.din0 (din_1_10),
	.din0_valid (din_valid_1_10),
	.din1 (din_1_11),
	.din1_valid (din_valid_1_11),
	.dout0 (dout_1_10),
	.dout0_valid (dout_valid_1_10),
	.dout1 (dout_1_11),
	.dout1_valid (dout_valid_1_11)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_6 (
	.clk (clk),
	.din0 (din_1_12),
	.din0_valid (din_valid_1_12),
	.din1 (din_1_13),
	.din1_valid (din_valid_1_13),
	.dout0 (dout_1_12),
	.dout0_valid (dout_valid_1_12),
	.dout1 (dout_1_13),
	.dout1_valid (dout_valid_1_13)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_7 (
	.clk (clk),
	.din0 (din_1_14),
	.din0_valid (din_valid_1_14),
	.din1 (din_1_15),
	.din1_valid (din_valid_1_15),
	.dout0 (dout_1_14),
	.dout0_valid (dout_valid_1_14),
	.dout1 (dout_1_15),
	.dout1_valid (dout_valid_1_15)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_8 (
	.clk (clk),
	.din0 (din_1_16),
	.din0_valid (din_valid_1_16),
	.din1 (din_1_17),
	.din1_valid (din_valid_1_17),
	.dout0 (dout_1_16),
	.dout0_valid (dout_valid_1_16),
	.dout1 (dout_1_17),
	.dout1_valid (dout_valid_1_17)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_9 (
	.clk (clk),
	.din0 (din_1_18),
	.din0_valid (din_valid_1_18),
	.din1 (din_1_19),
	.din1_valid (din_valid_1_19),
	.dout0 (dout_1_18),
	.dout0_valid (dout_valid_1_18),
	.dout1 (dout_1_19),
	.dout1_valid (dout_valid_1_19)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_10 (
	.clk (clk),
	.din0 (din_1_20),
	.din0_valid (din_valid_1_20),
	.din1 (din_1_21),
	.din1_valid (din_valid_1_21),
	.dout0 (dout_1_20),
	.dout0_valid (dout_valid_1_20),
	.dout1 (dout_1_21),
	.dout1_valid (dout_valid_1_21)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_11 (
	.clk (clk),
	.din0 (din_1_22),
	.din0_valid (din_valid_1_22),
	.din1 (din_1_23),
	.din1_valid (din_valid_1_23),
	.dout0 (dout_1_22),
	.dout0_valid (dout_valid_1_22),
	.dout1 (dout_1_23),
	.dout1_valid (dout_valid_1_23)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_12 (
	.clk (clk),
	.din0 (din_1_24),
	.din0_valid (din_valid_1_24),
	.din1 (din_1_25),
	.din1_valid (din_valid_1_25),
	.dout0 (dout_1_24),
	.dout0_valid (dout_valid_1_24),
	.dout1 (dout_1_25),
	.dout1_valid (dout_valid_1_25)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_13 (
	.clk (clk),
	.din0 (din_1_26),
	.din0_valid (din_valid_1_26),
	.din1 (din_1_27),
	.din1_valid (din_valid_1_27),
	.dout0 (dout_1_26),
	.dout0_valid (dout_valid_1_26),
	.dout1 (dout_1_27),
	.dout1_valid (dout_valid_1_27)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_14 (
	.clk (clk),
	.din0 (din_1_28),
	.din0_valid (din_valid_1_28),
	.din1 (din_1_29),
	.din1_valid (din_valid_1_29),
	.dout0 (dout_1_28),
	.dout0_valid (dout_valid_1_28),
	.dout1 (dout_1_29),
	.dout1_valid (dout_valid_1_29)
);

hashtable #(
	.ANDMSK(64'hffffffffffffffff),
	.NBITS(15),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(4096),
	.INIT_FILE("./mspm/string_matcher/bitmap1.mif")
)
hashtable_1_15 (
	.clk (clk),
	.din0 (din_1_30),
	.din0_valid (din_valid_1_30),
	.din1 (din_1_31),
	.din1_valid (din_valid_1_31),
	.dout0 (dout_1_30),
	.dout0_valid (dout_valid_1_30),
	.dout1 (dout_1_31),
	.dout1_valid (dout_valid_1_31)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_0 (
	.clk (clk),
	.din0 (din_2_0),
	.din0_valid (din_valid_2_0),
	.din1 (din_2_1),
	.din1_valid (din_valid_2_1),
	.dout0 (dout_2_0),
	.dout0_valid (dout_valid_2_0),
	.dout1 (dout_2_1),
	.dout1_valid (dout_valid_2_1)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_1 (
	.clk (clk),
	.din0 (din_2_2),
	.din0_valid (din_valid_2_2),
	.din1 (din_2_3),
	.din1_valid (din_valid_2_3),
	.dout0 (dout_2_2),
	.dout0_valid (dout_valid_2_2),
	.dout1 (dout_2_3),
	.dout1_valid (dout_valid_2_3)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_2 (
	.clk (clk),
	.din0 (din_2_4),
	.din0_valid (din_valid_2_4),
	.din1 (din_2_5),
	.din1_valid (din_valid_2_5),
	.dout0 (dout_2_4),
	.dout0_valid (dout_valid_2_4),
	.dout1 (dout_2_5),
	.dout1_valid (dout_valid_2_5)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_3 (
	.clk (clk),
	.din0 (din_2_6),
	.din0_valid (din_valid_2_6),
	.din1 (din_2_7),
	.din1_valid (din_valid_2_7),
	.dout0 (dout_2_6),
	.dout0_valid (dout_valid_2_6),
	.dout1 (dout_2_7),
	.dout1_valid (dout_valid_2_7)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_4 (
	.clk (clk),
	.din0 (din_2_8),
	.din0_valid (din_valid_2_8),
	.din1 (din_2_9),
	.din1_valid (din_valid_2_9),
	.dout0 (dout_2_8),
	.dout0_valid (dout_valid_2_8),
	.dout1 (dout_2_9),
	.dout1_valid (dout_valid_2_9)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_5 (
	.clk (clk),
	.din0 (din_2_10),
	.din0_valid (din_valid_2_10),
	.din1 (din_2_11),
	.din1_valid (din_valid_2_11),
	.dout0 (dout_2_10),
	.dout0_valid (dout_valid_2_10),
	.dout1 (dout_2_11),
	.dout1_valid (dout_valid_2_11)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_6 (
	.clk (clk),
	.din0 (din_2_12),
	.din0_valid (din_valid_2_12),
	.din1 (din_2_13),
	.din1_valid (din_valid_2_13),
	.dout0 (dout_2_12),
	.dout0_valid (dout_valid_2_12),
	.dout1 (dout_2_13),
	.dout1_valid (dout_valid_2_13)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_7 (
	.clk (clk),
	.din0 (din_2_14),
	.din0_valid (din_valid_2_14),
	.din1 (din_2_15),
	.din1_valid (din_valid_2_15),
	.dout0 (dout_2_14),
	.dout0_valid (dout_valid_2_14),
	.dout1 (dout_2_15),
	.dout1_valid (dout_valid_2_15)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_8 (
	.clk (clk),
	.din0 (din_2_16),
	.din0_valid (din_valid_2_16),
	.din1 (din_2_17),
	.din1_valid (din_valid_2_17),
	.dout0 (dout_2_16),
	.dout0_valid (dout_valid_2_16),
	.dout1 (dout_2_17),
	.dout1_valid (dout_valid_2_17)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_9 (
	.clk (clk),
	.din0 (din_2_18),
	.din0_valid (din_valid_2_18),
	.din1 (din_2_19),
	.din1_valid (din_valid_2_19),
	.dout0 (dout_2_18),
	.dout0_valid (dout_valid_2_18),
	.dout1 (dout_2_19),
	.dout1_valid (dout_valid_2_19)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_10 (
	.clk (clk),
	.din0 (din_2_20),
	.din0_valid (din_valid_2_20),
	.din1 (din_2_21),
	.din1_valid (din_valid_2_21),
	.dout0 (dout_2_20),
	.dout0_valid (dout_valid_2_20),
	.dout1 (dout_2_21),
	.dout1_valid (dout_valid_2_21)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_11 (
	.clk (clk),
	.din0 (din_2_22),
	.din0_valid (din_valid_2_22),
	.din1 (din_2_23),
	.din1_valid (din_valid_2_23),
	.dout0 (dout_2_22),
	.dout0_valid (dout_valid_2_22),
	.dout1 (dout_2_23),
	.dout1_valid (dout_valid_2_23)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_12 (
	.clk (clk),
	.din0 (din_2_24),
	.din0_valid (din_valid_2_24),
	.din1 (din_2_25),
	.din1_valid (din_valid_2_25),
	.dout0 (dout_2_24),
	.dout0_valid (dout_valid_2_24),
	.dout1 (dout_2_25),
	.dout1_valid (dout_valid_2_25)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_13 (
	.clk (clk),
	.din0 (din_2_26),
	.din0_valid (din_valid_2_26),
	.din1 (din_2_27),
	.din1_valid (din_valid_2_27),
	.dout0 (dout_2_26),
	.dout0_valid (dout_valid_2_26),
	.dout1 (dout_2_27),
	.dout1_valid (dout_valid_2_27)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_14 (
	.clk (clk),
	.din0 (din_2_28),
	.din0_valid (din_valid_2_28),
	.din1 (din_2_29),
	.din1_valid (din_valid_2_29),
	.dout0 (dout_2_28),
	.dout0_valid (dout_valid_2_28),
	.dout1 (dout_2_29),
	.dout1_valid (dout_valid_2_29)
);

hashtable #(
	.ANDMSK(64'hffffffffffffff00),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap2.mif")
)
hashtable_2_15 (
	.clk (clk),
	.din0 (din_2_30),
	.din0_valid (din_valid_2_30),
	.din1 (din_2_31),
	.din1_valid (din_valid_2_31),
	.dout0 (dout_2_30),
	.dout0_valid (dout_valid_2_30),
	.dout1 (dout_2_31),
	.dout1_valid (dout_valid_2_31)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_0 (
	.clk (clk),
	.din0 (din_3_0),
	.din0_valid (din_valid_3_0),
	.din1 (din_3_1),
	.din1_valid (din_valid_3_1),
	.dout0 (dout_3_0),
	.dout0_valid (dout_valid_3_0),
	.dout1 (dout_3_1),
	.dout1_valid (dout_valid_3_1)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_1 (
	.clk (clk),
	.din0 (din_3_2),
	.din0_valid (din_valid_3_2),
	.din1 (din_3_3),
	.din1_valid (din_valid_3_3),
	.dout0 (dout_3_2),
	.dout0_valid (dout_valid_3_2),
	.dout1 (dout_3_3),
	.dout1_valid (dout_valid_3_3)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_2 (
	.clk (clk),
	.din0 (din_3_4),
	.din0_valid (din_valid_3_4),
	.din1 (din_3_5),
	.din1_valid (din_valid_3_5),
	.dout0 (dout_3_4),
	.dout0_valid (dout_valid_3_4),
	.dout1 (dout_3_5),
	.dout1_valid (dout_valid_3_5)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_3 (
	.clk (clk),
	.din0 (din_3_6),
	.din0_valid (din_valid_3_6),
	.din1 (din_3_7),
	.din1_valid (din_valid_3_7),
	.dout0 (dout_3_6),
	.dout0_valid (dout_valid_3_6),
	.dout1 (dout_3_7),
	.dout1_valid (dout_valid_3_7)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_4 (
	.clk (clk),
	.din0 (din_3_8),
	.din0_valid (din_valid_3_8),
	.din1 (din_3_9),
	.din1_valid (din_valid_3_9),
	.dout0 (dout_3_8),
	.dout0_valid (dout_valid_3_8),
	.dout1 (dout_3_9),
	.dout1_valid (dout_valid_3_9)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_5 (
	.clk (clk),
	.din0 (din_3_10),
	.din0_valid (din_valid_3_10),
	.din1 (din_3_11),
	.din1_valid (din_valid_3_11),
	.dout0 (dout_3_10),
	.dout0_valid (dout_valid_3_10),
	.dout1 (dout_3_11),
	.dout1_valid (dout_valid_3_11)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_6 (
	.clk (clk),
	.din0 (din_3_12),
	.din0_valid (din_valid_3_12),
	.din1 (din_3_13),
	.din1_valid (din_valid_3_13),
	.dout0 (dout_3_12),
	.dout0_valid (dout_valid_3_12),
	.dout1 (dout_3_13),
	.dout1_valid (dout_valid_3_13)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_7 (
	.clk (clk),
	.din0 (din_3_14),
	.din0_valid (din_valid_3_14),
	.din1 (din_3_15),
	.din1_valid (din_valid_3_15),
	.dout0 (dout_3_14),
	.dout0_valid (dout_valid_3_14),
	.dout1 (dout_3_15),
	.dout1_valid (dout_valid_3_15)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_8 (
	.clk (clk),
	.din0 (din_3_16),
	.din0_valid (din_valid_3_16),
	.din1 (din_3_17),
	.din1_valid (din_valid_3_17),
	.dout0 (dout_3_16),
	.dout0_valid (dout_valid_3_16),
	.dout1 (dout_3_17),
	.dout1_valid (dout_valid_3_17)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_9 (
	.clk (clk),
	.din0 (din_3_18),
	.din0_valid (din_valid_3_18),
	.din1 (din_3_19),
	.din1_valid (din_valid_3_19),
	.dout0 (dout_3_18),
	.dout0_valid (dout_valid_3_18),
	.dout1 (dout_3_19),
	.dout1_valid (dout_valid_3_19)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_10 (
	.clk (clk),
	.din0 (din_3_20),
	.din0_valid (din_valid_3_20),
	.din1 (din_3_21),
	.din1_valid (din_valid_3_21),
	.dout0 (dout_3_20),
	.dout0_valid (dout_valid_3_20),
	.dout1 (dout_3_21),
	.dout1_valid (dout_valid_3_21)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_11 (
	.clk (clk),
	.din0 (din_3_22),
	.din0_valid (din_valid_3_22),
	.din1 (din_3_23),
	.din1_valid (din_valid_3_23),
	.dout0 (dout_3_22),
	.dout0_valid (dout_valid_3_22),
	.dout1 (dout_3_23),
	.dout1_valid (dout_valid_3_23)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_12 (
	.clk (clk),
	.din0 (din_3_24),
	.din0_valid (din_valid_3_24),
	.din1 (din_3_25),
	.din1_valid (din_valid_3_25),
	.dout0 (dout_3_24),
	.dout0_valid (dout_valid_3_24),
	.dout1 (dout_3_25),
	.dout1_valid (dout_valid_3_25)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_13 (
	.clk (clk),
	.din0 (din_3_26),
	.din0_valid (din_valid_3_26),
	.din1 (din_3_27),
	.din1_valid (din_valid_3_27),
	.dout0 (dout_3_26),
	.dout0_valid (dout_valid_3_26),
	.dout1 (dout_3_27),
	.dout1_valid (dout_valid_3_27)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_14 (
	.clk (clk),
	.din0 (din_3_28),
	.din0_valid (din_valid_3_28),
	.din1 (din_3_29),
	.din1_valid (din_valid_3_29),
	.dout0 (dout_3_28),
	.dout0_valid (dout_valid_3_28),
	.dout1 (dout_3_29),
	.dout1_valid (dout_valid_3_29)
);

hashtable #(
	.ANDMSK(64'hffffffffffff0000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap3.mif")
)
hashtable_3_15 (
	.clk (clk),
	.din0 (din_3_30),
	.din0_valid (din_valid_3_30),
	.din1 (din_3_31),
	.din1_valid (din_valid_3_31),
	.dout0 (dout_3_30),
	.dout0_valid (dout_valid_3_30),
	.dout1 (dout_3_31),
	.dout1_valid (dout_valid_3_31)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_0 (
	.clk (clk),
	.din0 (din_4_0),
	.din0_valid (din_valid_4_0),
	.din1 (din_4_1),
	.din1_valid (din_valid_4_1),
	.dout0 (dout_4_0),
	.dout0_valid (dout_valid_4_0),
	.dout1 (dout_4_1),
	.dout1_valid (dout_valid_4_1)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_1 (
	.clk (clk),
	.din0 (din_4_2),
	.din0_valid (din_valid_4_2),
	.din1 (din_4_3),
	.din1_valid (din_valid_4_3),
	.dout0 (dout_4_2),
	.dout0_valid (dout_valid_4_2),
	.dout1 (dout_4_3),
	.dout1_valid (dout_valid_4_3)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_2 (
	.clk (clk),
	.din0 (din_4_4),
	.din0_valid (din_valid_4_4),
	.din1 (din_4_5),
	.din1_valid (din_valid_4_5),
	.dout0 (dout_4_4),
	.dout0_valid (dout_valid_4_4),
	.dout1 (dout_4_5),
	.dout1_valid (dout_valid_4_5)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_3 (
	.clk (clk),
	.din0 (din_4_6),
	.din0_valid (din_valid_4_6),
	.din1 (din_4_7),
	.din1_valid (din_valid_4_7),
	.dout0 (dout_4_6),
	.dout0_valid (dout_valid_4_6),
	.dout1 (dout_4_7),
	.dout1_valid (dout_valid_4_7)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_4 (
	.clk (clk),
	.din0 (din_4_8),
	.din0_valid (din_valid_4_8),
	.din1 (din_4_9),
	.din1_valid (din_valid_4_9),
	.dout0 (dout_4_8),
	.dout0_valid (dout_valid_4_8),
	.dout1 (dout_4_9),
	.dout1_valid (dout_valid_4_9)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_5 (
	.clk (clk),
	.din0 (din_4_10),
	.din0_valid (din_valid_4_10),
	.din1 (din_4_11),
	.din1_valid (din_valid_4_11),
	.dout0 (dout_4_10),
	.dout0_valid (dout_valid_4_10),
	.dout1 (dout_4_11),
	.dout1_valid (dout_valid_4_11)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_6 (
	.clk (clk),
	.din0 (din_4_12),
	.din0_valid (din_valid_4_12),
	.din1 (din_4_13),
	.din1_valid (din_valid_4_13),
	.dout0 (dout_4_12),
	.dout0_valid (dout_valid_4_12),
	.dout1 (dout_4_13),
	.dout1_valid (dout_valid_4_13)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_7 (
	.clk (clk),
	.din0 (din_4_14),
	.din0_valid (din_valid_4_14),
	.din1 (din_4_15),
	.din1_valid (din_valid_4_15),
	.dout0 (dout_4_14),
	.dout0_valid (dout_valid_4_14),
	.dout1 (dout_4_15),
	.dout1_valid (dout_valid_4_15)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_8 (
	.clk (clk),
	.din0 (din_4_16),
	.din0_valid (din_valid_4_16),
	.din1 (din_4_17),
	.din1_valid (din_valid_4_17),
	.dout0 (dout_4_16),
	.dout0_valid (dout_valid_4_16),
	.dout1 (dout_4_17),
	.dout1_valid (dout_valid_4_17)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_9 (
	.clk (clk),
	.din0 (din_4_18),
	.din0_valid (din_valid_4_18),
	.din1 (din_4_19),
	.din1_valid (din_valid_4_19),
	.dout0 (dout_4_18),
	.dout0_valid (dout_valid_4_18),
	.dout1 (dout_4_19),
	.dout1_valid (dout_valid_4_19)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_10 (
	.clk (clk),
	.din0 (din_4_20),
	.din0_valid (din_valid_4_20),
	.din1 (din_4_21),
	.din1_valid (din_valid_4_21),
	.dout0 (dout_4_20),
	.dout0_valid (dout_valid_4_20),
	.dout1 (dout_4_21),
	.dout1_valid (dout_valid_4_21)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_11 (
	.clk (clk),
	.din0 (din_4_22),
	.din0_valid (din_valid_4_22),
	.din1 (din_4_23),
	.din1_valid (din_valid_4_23),
	.dout0 (dout_4_22),
	.dout0_valid (dout_valid_4_22),
	.dout1 (dout_4_23),
	.dout1_valid (dout_valid_4_23)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_12 (
	.clk (clk),
	.din0 (din_4_24),
	.din0_valid (din_valid_4_24),
	.din1 (din_4_25),
	.din1_valid (din_valid_4_25),
	.dout0 (dout_4_24),
	.dout0_valid (dout_valid_4_24),
	.dout1 (dout_4_25),
	.dout1_valid (dout_valid_4_25)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_13 (
	.clk (clk),
	.din0 (din_4_26),
	.din0_valid (din_valid_4_26),
	.din1 (din_4_27),
	.din1_valid (din_valid_4_27),
	.dout0 (dout_4_26),
	.dout0_valid (dout_valid_4_26),
	.dout1 (dout_4_27),
	.dout1_valid (dout_valid_4_27)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_14 (
	.clk (clk),
	.din0 (din_4_28),
	.din0_valid (din_valid_4_28),
	.din1 (din_4_29),
	.din1_valid (din_valid_4_29),
	.dout0 (dout_4_28),
	.dout0_valid (dout_valid_4_28),
	.dout1 (dout_4_29),
	.dout1_valid (dout_valid_4_29)
);

hashtable #(
	.ANDMSK(64'hffffffffff000000),
	.NBITS(11),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(256),
	.INIT_FILE("./mspm/string_matcher/bitmap4.mif")
)
hashtable_4_15 (
	.clk (clk),
	.din0 (din_4_30),
	.din0_valid (din_valid_4_30),
	.din1 (din_4_31),
	.din1_valid (din_valid_4_31),
	.dout0 (dout_4_30),
	.dout0_valid (dout_valid_4_30),
	.dout1 (dout_4_31),
	.dout1_valid (dout_valid_4_31)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_0 (
	.clk (clk),
	.din0 (din_5_0),
	.din0_valid (din_valid_5_0),
	.din1 (din_5_1),
	.din1_valid (din_valid_5_1),
	.dout0 (dout_5_0),
	.dout0_valid (dout_valid_5_0),
	.dout1 (dout_5_1),
	.dout1_valid (dout_valid_5_1)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_1 (
	.clk (clk),
	.din0 (din_5_2),
	.din0_valid (din_valid_5_2),
	.din1 (din_5_3),
	.din1_valid (din_valid_5_3),
	.dout0 (dout_5_2),
	.dout0_valid (dout_valid_5_2),
	.dout1 (dout_5_3),
	.dout1_valid (dout_valid_5_3)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_2 (
	.clk (clk),
	.din0 (din_5_4),
	.din0_valid (din_valid_5_4),
	.din1 (din_5_5),
	.din1_valid (din_valid_5_5),
	.dout0 (dout_5_4),
	.dout0_valid (dout_valid_5_4),
	.dout1 (dout_5_5),
	.dout1_valid (dout_valid_5_5)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_3 (
	.clk (clk),
	.din0 (din_5_6),
	.din0_valid (din_valid_5_6),
	.din1 (din_5_7),
	.din1_valid (din_valid_5_7),
	.dout0 (dout_5_6),
	.dout0_valid (dout_valid_5_6),
	.dout1 (dout_5_7),
	.dout1_valid (dout_valid_5_7)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_4 (
	.clk (clk),
	.din0 (din_5_8),
	.din0_valid (din_valid_5_8),
	.din1 (din_5_9),
	.din1_valid (din_valid_5_9),
	.dout0 (dout_5_8),
	.dout0_valid (dout_valid_5_8),
	.dout1 (dout_5_9),
	.dout1_valid (dout_valid_5_9)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_5 (
	.clk (clk),
	.din0 (din_5_10),
	.din0_valid (din_valid_5_10),
	.din1 (din_5_11),
	.din1_valid (din_valid_5_11),
	.dout0 (dout_5_10),
	.dout0_valid (dout_valid_5_10),
	.dout1 (dout_5_11),
	.dout1_valid (dout_valid_5_11)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_6 (
	.clk (clk),
	.din0 (din_5_12),
	.din0_valid (din_valid_5_12),
	.din1 (din_5_13),
	.din1_valid (din_valid_5_13),
	.dout0 (dout_5_12),
	.dout0_valid (dout_valid_5_12),
	.dout1 (dout_5_13),
	.dout1_valid (dout_valid_5_13)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_7 (
	.clk (clk),
	.din0 (din_5_14),
	.din0_valid (din_valid_5_14),
	.din1 (din_5_15),
	.din1_valid (din_valid_5_15),
	.dout0 (dout_5_14),
	.dout0_valid (dout_valid_5_14),
	.dout1 (dout_5_15),
	.dout1_valid (dout_valid_5_15)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_8 (
	.clk (clk),
	.din0 (din_5_16),
	.din0_valid (din_valid_5_16),
	.din1 (din_5_17),
	.din1_valid (din_valid_5_17),
	.dout0 (dout_5_16),
	.dout0_valid (dout_valid_5_16),
	.dout1 (dout_5_17),
	.dout1_valid (dout_valid_5_17)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_9 (
	.clk (clk),
	.din0 (din_5_18),
	.din0_valid (din_valid_5_18),
	.din1 (din_5_19),
	.din1_valid (din_valid_5_19),
	.dout0 (dout_5_18),
	.dout0_valid (dout_valid_5_18),
	.dout1 (dout_5_19),
	.dout1_valid (dout_valid_5_19)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_10 (
	.clk (clk),
	.din0 (din_5_20),
	.din0_valid (din_valid_5_20),
	.din1 (din_5_21),
	.din1_valid (din_valid_5_21),
	.dout0 (dout_5_20),
	.dout0_valid (dout_valid_5_20),
	.dout1 (dout_5_21),
	.dout1_valid (dout_valid_5_21)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_11 (
	.clk (clk),
	.din0 (din_5_22),
	.din0_valid (din_valid_5_22),
	.din1 (din_5_23),
	.din1_valid (din_valid_5_23),
	.dout0 (dout_5_22),
	.dout0_valid (dout_valid_5_22),
	.dout1 (dout_5_23),
	.dout1_valid (dout_valid_5_23)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_12 (
	.clk (clk),
	.din0 (din_5_24),
	.din0_valid (din_valid_5_24),
	.din1 (din_5_25),
	.din1_valid (din_valid_5_25),
	.dout0 (dout_5_24),
	.dout0_valid (dout_valid_5_24),
	.dout1 (dout_5_25),
	.dout1_valid (dout_valid_5_25)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_13 (
	.clk (clk),
	.din0 (din_5_26),
	.din0_valid (din_valid_5_26),
	.din1 (din_5_27),
	.din1_valid (din_valid_5_27),
	.dout0 (dout_5_26),
	.dout0_valid (dout_valid_5_26),
	.dout1 (dout_5_27),
	.dout1_valid (dout_valid_5_27)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_14 (
	.clk (clk),
	.din0 (din_5_28),
	.din0_valid (din_valid_5_28),
	.din1 (din_5_29),
	.din1_valid (din_valid_5_29),
	.dout0 (dout_5_28),
	.dout0_valid (dout_valid_5_28),
	.dout1 (dout_5_29),
	.dout1_valid (dout_valid_5_29)
);

hashtable #(
	.ANDMSK(64'hffffffff00000000),
	.NBITS(12),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(512),
	.INIT_FILE("./mspm/string_matcher/bitmap5.mif")
)
hashtable_5_15 (
	.clk (clk),
	.din0 (din_5_30),
	.din0_valid (din_valid_5_30),
	.din1 (din_5_31),
	.din1_valid (din_valid_5_31),
	.dout0 (dout_5_30),
	.dout0_valid (dout_valid_5_30),
	.dout1 (dout_5_31),
	.dout1_valid (dout_valid_5_31)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_0 (
	.clk (clk),
	.din0 (din_6_0),
	.din0_valid (din_valid_6_0),
	.din1 (din_6_1),
	.din1_valid (din_valid_6_1),
	.dout0 (dout_6_0),
	.dout0_valid (dout_valid_6_0),
	.dout1 (dout_6_1),
	.dout1_valid (dout_valid_6_1)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_1 (
	.clk (clk),
	.din0 (din_6_2),
	.din0_valid (din_valid_6_2),
	.din1 (din_6_3),
	.din1_valid (din_valid_6_3),
	.dout0 (dout_6_2),
	.dout0_valid (dout_valid_6_2),
	.dout1 (dout_6_3),
	.dout1_valid (dout_valid_6_3)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_2 (
	.clk (clk),
	.din0 (din_6_4),
	.din0_valid (din_valid_6_4),
	.din1 (din_6_5),
	.din1_valid (din_valid_6_5),
	.dout0 (dout_6_4),
	.dout0_valid (dout_valid_6_4),
	.dout1 (dout_6_5),
	.dout1_valid (dout_valid_6_5)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_3 (
	.clk (clk),
	.din0 (din_6_6),
	.din0_valid (din_valid_6_6),
	.din1 (din_6_7),
	.din1_valid (din_valid_6_7),
	.dout0 (dout_6_6),
	.dout0_valid (dout_valid_6_6),
	.dout1 (dout_6_7),
	.dout1_valid (dout_valid_6_7)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_4 (
	.clk (clk),
	.din0 (din_6_8),
	.din0_valid (din_valid_6_8),
	.din1 (din_6_9),
	.din1_valid (din_valid_6_9),
	.dout0 (dout_6_8),
	.dout0_valid (dout_valid_6_8),
	.dout1 (dout_6_9),
	.dout1_valid (dout_valid_6_9)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_5 (
	.clk (clk),
	.din0 (din_6_10),
	.din0_valid (din_valid_6_10),
	.din1 (din_6_11),
	.din1_valid (din_valid_6_11),
	.dout0 (dout_6_10),
	.dout0_valid (dout_valid_6_10),
	.dout1 (dout_6_11),
	.dout1_valid (dout_valid_6_11)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_6 (
	.clk (clk),
	.din0 (din_6_12),
	.din0_valid (din_valid_6_12),
	.din1 (din_6_13),
	.din1_valid (din_valid_6_13),
	.dout0 (dout_6_12),
	.dout0_valid (dout_valid_6_12),
	.dout1 (dout_6_13),
	.dout1_valid (dout_valid_6_13)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_7 (
	.clk (clk),
	.din0 (din_6_14),
	.din0_valid (din_valid_6_14),
	.din1 (din_6_15),
	.din1_valid (din_valid_6_15),
	.dout0 (dout_6_14),
	.dout0_valid (dout_valid_6_14),
	.dout1 (dout_6_15),
	.dout1_valid (dout_valid_6_15)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_8 (
	.clk (clk),
	.din0 (din_6_16),
	.din0_valid (din_valid_6_16),
	.din1 (din_6_17),
	.din1_valid (din_valid_6_17),
	.dout0 (dout_6_16),
	.dout0_valid (dout_valid_6_16),
	.dout1 (dout_6_17),
	.dout1_valid (dout_valid_6_17)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_9 (
	.clk (clk),
	.din0 (din_6_18),
	.din0_valid (din_valid_6_18),
	.din1 (din_6_19),
	.din1_valid (din_valid_6_19),
	.dout0 (dout_6_18),
	.dout0_valid (dout_valid_6_18),
	.dout1 (dout_6_19),
	.dout1_valid (dout_valid_6_19)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_10 (
	.clk (clk),
	.din0 (din_6_20),
	.din0_valid (din_valid_6_20),
	.din1 (din_6_21),
	.din1_valid (din_valid_6_21),
	.dout0 (dout_6_20),
	.dout0_valid (dout_valid_6_20),
	.dout1 (dout_6_21),
	.dout1_valid (dout_valid_6_21)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_11 (
	.clk (clk),
	.din0 (din_6_22),
	.din0_valid (din_valid_6_22),
	.din1 (din_6_23),
	.din1_valid (din_valid_6_23),
	.dout0 (dout_6_22),
	.dout0_valid (dout_valid_6_22),
	.dout1 (dout_6_23),
	.dout1_valid (dout_valid_6_23)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_12 (
	.clk (clk),
	.din0 (din_6_24),
	.din0_valid (din_valid_6_24),
	.din1 (din_6_25),
	.din1_valid (din_valid_6_25),
	.dout0 (dout_6_24),
	.dout0_valid (dout_valid_6_24),
	.dout1 (dout_6_25),
	.dout1_valid (dout_valid_6_25)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_13 (
	.clk (clk),
	.din0 (din_6_26),
	.din0_valid (din_valid_6_26),
	.din1 (din_6_27),
	.din1_valid (din_valid_6_27),
	.dout0 (dout_6_26),
	.dout0_valid (dout_valid_6_26),
	.dout1 (dout_6_27),
	.dout1_valid (dout_valid_6_27)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_14 (
	.clk (clk),
	.din0 (din_6_28),
	.din0_valid (din_valid_6_28),
	.din1 (din_6_29),
	.din1_valid (din_valid_6_29),
	.dout0 (dout_6_28),
	.dout0_valid (dout_valid_6_28),
	.dout1 (dout_6_29),
	.dout1_valid (dout_valid_6_29)
);

hashtable #(
	.ANDMSK(64'hffffff0000000000),
	.NBITS(10),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(128),
	.INIT_FILE("./mspm/string_matcher/bitmap6.mif")
)
hashtable_6_15 (
	.clk (clk),
	.din0 (din_6_30),
	.din0_valid (din_valid_6_30),
	.din1 (din_6_31),
	.din1_valid (din_valid_6_31),
	.dout0 (dout_6_30),
	.dout0_valid (dout_valid_6_30),
	.dout1 (dout_6_31),
	.dout1_valid (dout_valid_6_31)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_0 (
	.clk (clk),
	.din0 (din_7_0),
	.din0_valid (din_valid_7_0),
	.din1 (din_7_1),
	.din1_valid (din_valid_7_1),
	.dout0 (dout_7_0),
	.dout0_valid (dout_valid_7_0),
	.dout1 (dout_7_1),
	.dout1_valid (dout_valid_7_1)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_1 (
	.clk (clk),
	.din0 (din_7_2),
	.din0_valid (din_valid_7_2),
	.din1 (din_7_3),
	.din1_valid (din_valid_7_3),
	.dout0 (dout_7_2),
	.dout0_valid (dout_valid_7_2),
	.dout1 (dout_7_3),
	.dout1_valid (dout_valid_7_3)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_2 (
	.clk (clk),
	.din0 (din_7_4),
	.din0_valid (din_valid_7_4),
	.din1 (din_7_5),
	.din1_valid (din_valid_7_5),
	.dout0 (dout_7_4),
	.dout0_valid (dout_valid_7_4),
	.dout1 (dout_7_5),
	.dout1_valid (dout_valid_7_5)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_3 (
	.clk (clk),
	.din0 (din_7_6),
	.din0_valid (din_valid_7_6),
	.din1 (din_7_7),
	.din1_valid (din_valid_7_7),
	.dout0 (dout_7_6),
	.dout0_valid (dout_valid_7_6),
	.dout1 (dout_7_7),
	.dout1_valid (dout_valid_7_7)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_4 (
	.clk (clk),
	.din0 (din_7_8),
	.din0_valid (din_valid_7_8),
	.din1 (din_7_9),
	.din1_valid (din_valid_7_9),
	.dout0 (dout_7_8),
	.dout0_valid (dout_valid_7_8),
	.dout1 (dout_7_9),
	.dout1_valid (dout_valid_7_9)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_5 (
	.clk (clk),
	.din0 (din_7_10),
	.din0_valid (din_valid_7_10),
	.din1 (din_7_11),
	.din1_valid (din_valid_7_11),
	.dout0 (dout_7_10),
	.dout0_valid (dout_valid_7_10),
	.dout1 (dout_7_11),
	.dout1_valid (dout_valid_7_11)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_6 (
	.clk (clk),
	.din0 (din_7_12),
	.din0_valid (din_valid_7_12),
	.din1 (din_7_13),
	.din1_valid (din_valid_7_13),
	.dout0 (dout_7_12),
	.dout0_valid (dout_valid_7_12),
	.dout1 (dout_7_13),
	.dout1_valid (dout_valid_7_13)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_7 (
	.clk (clk),
	.din0 (din_7_14),
	.din0_valid (din_valid_7_14),
	.din1 (din_7_15),
	.din1_valid (din_valid_7_15),
	.dout0 (dout_7_14),
	.dout0_valid (dout_valid_7_14),
	.dout1 (dout_7_15),
	.dout1_valid (dout_valid_7_15)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_8 (
	.clk (clk),
	.din0 (din_7_16),
	.din0_valid (din_valid_7_16),
	.din1 (din_7_17),
	.din1_valid (din_valid_7_17),
	.dout0 (dout_7_16),
	.dout0_valid (dout_valid_7_16),
	.dout1 (dout_7_17),
	.dout1_valid (dout_valid_7_17)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_9 (
	.clk (clk),
	.din0 (din_7_18),
	.din0_valid (din_valid_7_18),
	.din1 (din_7_19),
	.din1_valid (din_valid_7_19),
	.dout0 (dout_7_18),
	.dout0_valid (dout_valid_7_18),
	.dout1 (dout_7_19),
	.dout1_valid (dout_valid_7_19)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_10 (
	.clk (clk),
	.din0 (din_7_20),
	.din0_valid (din_valid_7_20),
	.din1 (din_7_21),
	.din1_valid (din_valid_7_21),
	.dout0 (dout_7_20),
	.dout0_valid (dout_valid_7_20),
	.dout1 (dout_7_21),
	.dout1_valid (dout_valid_7_21)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_11 (
	.clk (clk),
	.din0 (din_7_22),
	.din0_valid (din_valid_7_22),
	.din1 (din_7_23),
	.din1_valid (din_valid_7_23),
	.dout0 (dout_7_22),
	.dout0_valid (dout_valid_7_22),
	.dout1 (dout_7_23),
	.dout1_valid (dout_valid_7_23)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_12 (
	.clk (clk),
	.din0 (din_7_24),
	.din0_valid (din_valid_7_24),
	.din1 (din_7_25),
	.din1_valid (din_valid_7_25),
	.dout0 (dout_7_24),
	.dout0_valid (dout_valid_7_24),
	.dout1 (dout_7_25),
	.dout1_valid (dout_valid_7_25)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_13 (
	.clk (clk),
	.din0 (din_7_26),
	.din0_valid (din_valid_7_26),
	.din1 (din_7_27),
	.din1_valid (din_valid_7_27),
	.dout0 (dout_7_26),
	.dout0_valid (dout_valid_7_26),
	.dout1 (dout_7_27),
	.dout1_valid (dout_valid_7_27)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_14 (
	.clk (clk),
	.din0 (din_7_28),
	.din0_valid (din_valid_7_28),
	.din1 (din_7_29),
	.din1_valid (din_valid_7_29),
	.dout0 (dout_7_28),
	.dout0_valid (dout_valid_7_28),
	.dout1 (dout_7_29),
	.dout1_valid (dout_valid_7_29)
);

hashtable #(
	.ANDMSK(64'hffff000000000000),
	.NBITS(8),
	.DWIDTH(RID_WIDTH),
	.MEM_SIZE(32),
	.INIT_FILE("./mspm/string_matcher/bitmap7.mif")
)
hashtable_7_15 (
	.clk (clk),
	.din0 (din_7_30),
	.din0_valid (din_valid_7_30),
	.din1 (din_7_31),
	.din1_valid (din_valid_7_31),
	.dout0 (dout_7_30),
	.dout0_valid (dout_valid_7_30),
	.dout1 (dout_7_31),
	.dout1_valid (dout_valid_7_31)
);

endmodule
